-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity initInputs is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    matrix_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    matrix_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    matrix_in_pipe_read_data : in   std_logic_vector(15 downto 0);
    maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initInputs;
architecture initInputs_arch of initInputs is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal initInputs_CP_117_start: Boolean;
  signal initInputs_CP_117_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_263_store_0_req_1 : boolean;
  signal ptr_deref_263_store_0_ack_1 : boolean;
  signal ptr_deref_259_store_0_ack_0 : boolean;
  signal ptr_deref_259_store_0_req_0 : boolean;
  signal ptr_deref_263_store_0_req_0 : boolean;
  signal ptr_deref_263_store_0_ack_0 : boolean;
  signal type_cast_233_inst_ack_1 : boolean;
  signal type_cast_233_inst_req_1 : boolean;
  signal ptr_deref_271_load_0_req_0 : boolean;
  signal ptr_deref_271_load_0_ack_0 : boolean;
  signal type_cast_233_inst_ack_0 : boolean;
  signal type_cast_233_inst_req_0 : boolean;
  signal ptr_deref_259_store_0_ack_1 : boolean;
  signal type_cast_256_inst_ack_1 : boolean;
  signal ptr_deref_259_store_0_req_1 : boolean;
  signal ptr_deref_243_load_0_ack_1 : boolean;
  signal ptr_deref_243_load_0_req_1 : boolean;
  signal ptr_deref_203_load_0_ack_1 : boolean;
  signal ptr_deref_229_load_0_ack_1 : boolean;
  signal ptr_deref_229_load_0_req_1 : boolean;
  signal ptr_deref_83_load_0_req_0 : boolean;
  signal ptr_deref_83_load_0_ack_0 : boolean;
  signal ptr_deref_83_load_0_req_1 : boolean;
  signal ptr_deref_83_load_0_ack_1 : boolean;
  signal ptr_deref_229_load_0_ack_0 : boolean;
  signal ptr_deref_229_load_0_req_0 : boolean;
  signal ptr_deref_203_load_0_req_1 : boolean;
  signal RPIPE_maxNitr_in_75_inst_req_0 : boolean;
  signal RPIPE_maxNitr_in_75_inst_ack_0 : boolean;
  signal RPIPE_maxNitr_in_75_inst_req_1 : boolean;
  signal RPIPE_maxNitr_in_75_inst_ack_1 : boolean;
  signal ADD_u32_u32_252_inst_ack_0 : boolean;
  signal ADD_u32_u32_252_inst_req_0 : boolean;
  signal type_cast_256_inst_req_1 : boolean;
  signal ptr_deref_78_store_0_req_0 : boolean;
  signal ptr_deref_78_store_0_ack_0 : boolean;
  signal ptr_deref_78_store_0_req_1 : boolean;
  signal ptr_deref_78_store_0_ack_1 : boolean;
  signal type_cast_247_inst_ack_1 : boolean;
  signal type_cast_247_inst_req_1 : boolean;
  signal type_cast_247_inst_ack_0 : boolean;
  signal STORE_ncol_ind_218_store_0_ack_1 : boolean;
  signal STORE_ncol_ind_218_store_0_req_1 : boolean;
  signal STORE_maxNitr_85_store_0_req_0 : boolean;
  signal STORE_maxNitr_85_store_0_ack_0 : boolean;
  signal STORE_maxNitr_85_store_0_req_1 : boolean;
  signal STORE_maxNitr_85_store_0_ack_1 : boolean;
  signal type_cast_247_inst_req_0 : boolean;
  signal RPIPE_ebbyNo_in_89_inst_req_0 : boolean;
  signal RPIPE_ebbyNo_in_89_inst_ack_0 : boolean;
  signal STORE_ncol_ind_218_store_0_ack_0 : boolean;
  signal RPIPE_ebbyNo_in_89_inst_req_1 : boolean;
  signal RPIPE_ebbyNo_in_89_inst_ack_1 : boolean;
  signal ADD_u32_u32_252_inst_ack_1 : boolean;
  signal STORE_ncol_ind_218_store_0_req_0 : boolean;
  signal ptr_deref_92_store_0_req_0 : boolean;
  signal ptr_deref_92_store_0_ack_0 : boolean;
  signal ptr_deref_92_store_0_req_1 : boolean;
  signal ptr_deref_92_store_0_ack_1 : boolean;
  signal ptr_deref_243_load_0_ack_0 : boolean;
  signal ptr_deref_243_load_0_req_0 : boolean;
  signal ptr_deref_97_load_0_req_0 : boolean;
  signal ptr_deref_97_load_0_ack_0 : boolean;
  signal ptr_deref_97_load_0_req_1 : boolean;
  signal ptr_deref_97_load_0_ack_1 : boolean;
  signal ptr_deref_216_load_0_ack_1 : boolean;
  signal ptr_deref_216_load_0_req_1 : boolean;
  signal STORE_ebbyNo_99_store_0_req_0 : boolean;
  signal STORE_ebbyNo_99_store_0_ack_0 : boolean;
  signal STORE_ebbyNo_99_store_0_req_1 : boolean;
  signal STORE_ebbyNo_99_store_0_ack_1 : boolean;
  signal type_cast_256_inst_ack_0 : boolean;
  signal ptr_deref_216_load_0_ack_0 : boolean;
  signal ptr_deref_216_load_0_req_0 : boolean;
  signal ptr_deref_103_store_0_req_0 : boolean;
  signal ptr_deref_103_store_0_ack_0 : boolean;
  signal ptr_deref_103_store_0_req_1 : boolean;
  signal ptr_deref_103_store_0_ack_1 : boolean;
  signal ptr_deref_203_load_0_ack_0 : boolean;
  signal ptr_deref_111_load_0_req_0 : boolean;
  signal ptr_deref_111_load_0_ack_0 : boolean;
  signal ptr_deref_111_load_0_req_1 : boolean;
  signal ptr_deref_111_load_0_ack_1 : boolean;
  signal ptr_deref_203_load_0_req_0 : boolean;
  signal type_cast_116_inst_req_0 : boolean;
  signal type_cast_116_inst_ack_0 : boolean;
  signal type_cast_116_inst_req_1 : boolean;
  signal type_cast_116_inst_ack_1 : boolean;
  signal SLT_i32_u1_125_inst_req_0 : boolean;
  signal SLT_i32_u1_125_inst_ack_0 : boolean;
  signal SLT_i32_u1_125_inst_req_1 : boolean;
  signal SLT_i32_u1_125_inst_ack_1 : boolean;
  signal type_cast_256_inst_req_0 : boolean;
  signal if_stmt_128_branch_req_0 : boolean;
  signal if_stmt_128_branch_ack_1 : boolean;
  signal if_stmt_128_branch_ack_0 : boolean;
  signal STORE_ncols_205_store_0_ack_1 : boolean;
  signal STORE_ncols_205_store_0_req_1 : boolean;
  signal RPIPE_matrix_in_136_inst_req_0 : boolean;
  signal RPIPE_matrix_in_136_inst_ack_0 : boolean;
  signal RPIPE_matrix_in_136_inst_req_1 : boolean;
  signal RPIPE_matrix_in_136_inst_ack_1 : boolean;
  signal ADD_u32_u32_252_inst_req_1 : boolean;
  signal STORE_ncols_205_store_0_ack_0 : boolean;
  signal STORE_ncols_205_store_0_req_0 : boolean;
  signal ptr_deref_139_store_0_req_0 : boolean;
  signal ptr_deref_139_store_0_ack_0 : boolean;
  signal ptr_deref_139_store_0_req_1 : boolean;
  signal ptr_deref_139_store_0_ack_1 : boolean;
  signal ptr_deref_144_load_0_req_0 : boolean;
  signal ptr_deref_144_load_0_ack_0 : boolean;
  signal ptr_deref_144_load_0_req_1 : boolean;
  signal ptr_deref_144_load_0_ack_1 : boolean;
  signal ptr_deref_148_load_0_req_0 : boolean;
  signal ptr_deref_148_load_0_ack_0 : boolean;
  signal ptr_deref_148_load_0_req_1 : boolean;
  signal ptr_deref_148_load_0_ack_1 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal addr_of_158_final_reg_req_0 : boolean;
  signal addr_of_158_final_reg_ack_0 : boolean;
  signal addr_of_158_final_reg_req_1 : boolean;
  signal addr_of_158_final_reg_ack_1 : boolean;
  signal ptr_deref_161_store_0_req_0 : boolean;
  signal ptr_deref_161_store_0_ack_0 : boolean;
  signal ptr_deref_161_store_0_req_1 : boolean;
  signal ptr_deref_161_store_0_ack_1 : boolean;
  signal ptr_deref_168_load_0_req_0 : boolean;
  signal ptr_deref_168_load_0_ack_0 : boolean;
  signal ptr_deref_168_load_0_req_1 : boolean;
  signal ptr_deref_168_load_0_ack_1 : boolean;
  signal ADD_u16_u16_174_inst_req_0 : boolean;
  signal ADD_u16_u16_174_inst_ack_0 : boolean;
  signal ADD_u16_u16_174_inst_req_1 : boolean;
  signal ADD_u16_u16_174_inst_ack_1 : boolean;
  signal ptr_deref_177_store_0_req_0 : boolean;
  signal ptr_deref_177_store_0_ack_0 : boolean;
  signal ptr_deref_177_store_0_req_1 : boolean;
  signal ptr_deref_177_store_0_ack_1 : boolean;
  signal ptr_deref_190_load_0_req_0 : boolean;
  signal ptr_deref_190_load_0_ack_0 : boolean;
  signal ptr_deref_190_load_0_req_1 : boolean;
  signal ptr_deref_190_load_0_ack_1 : boolean;
  signal STORE_nrows_192_store_0_req_0 : boolean;
  signal STORE_nrows_192_store_0_ack_0 : boolean;
  signal STORE_nrows_192_store_0_req_1 : boolean;
  signal STORE_nrows_192_store_0_ack_1 : boolean;
  signal ptr_deref_271_load_0_req_1 : boolean;
  signal ptr_deref_271_load_0_ack_1 : boolean;
  signal type_cast_275_inst_req_0 : boolean;
  signal type_cast_275_inst_ack_0 : boolean;
  signal type_cast_275_inst_req_1 : boolean;
  signal type_cast_275_inst_ack_1 : boolean;
  signal ptr_deref_279_load_0_req_0 : boolean;
  signal ptr_deref_279_load_0_ack_0 : boolean;
  signal ptr_deref_279_load_0_req_1 : boolean;
  signal ptr_deref_279_load_0_ack_1 : boolean;
  signal type_cast_283_inst_req_0 : boolean;
  signal type_cast_283_inst_ack_0 : boolean;
  signal type_cast_283_inst_req_1 : boolean;
  signal type_cast_283_inst_ack_1 : boolean;
  signal SLT_i32_u1_290_inst_req_0 : boolean;
  signal SLT_i32_u1_290_inst_ack_0 : boolean;
  signal SLT_i32_u1_290_inst_req_1 : boolean;
  signal SLT_i32_u1_290_inst_ack_1 : boolean;
  signal if_stmt_292_branch_req_0 : boolean;
  signal if_stmt_292_branch_ack_1 : boolean;
  signal if_stmt_292_branch_ack_0 : boolean;
  signal RPIPE_matrix_in_300_inst_req_0 : boolean;
  signal RPIPE_matrix_in_300_inst_ack_0 : boolean;
  signal RPIPE_matrix_in_300_inst_req_1 : boolean;
  signal RPIPE_matrix_in_300_inst_ack_1 : boolean;
  signal ptr_deref_303_store_0_req_0 : boolean;
  signal ptr_deref_303_store_0_ack_0 : boolean;
  signal ptr_deref_303_store_0_req_1 : boolean;
  signal ptr_deref_303_store_0_ack_1 : boolean;
  signal ptr_deref_308_load_0_req_0 : boolean;
  signal ptr_deref_308_load_0_ack_0 : boolean;
  signal ptr_deref_308_load_0_req_1 : boolean;
  signal ptr_deref_308_load_0_ack_1 : boolean;
  signal ptr_deref_312_load_0_req_0 : boolean;
  signal ptr_deref_312_load_0_ack_0 : boolean;
  signal ptr_deref_312_load_0_req_1 : boolean;
  signal ptr_deref_312_load_0_ack_1 : boolean;
  signal type_cast_316_inst_req_0 : boolean;
  signal type_cast_316_inst_ack_0 : boolean;
  signal type_cast_316_inst_req_1 : boolean;
  signal type_cast_316_inst_ack_1 : boolean;
  signal ADD_u32_u32_322_inst_req_0 : boolean;
  signal ADD_u32_u32_322_inst_ack_0 : boolean;
  signal ADD_u32_u32_322_inst_req_1 : boolean;
  signal ADD_u32_u32_322_inst_ack_1 : boolean;
  signal type_cast_327_inst_req_0 : boolean;
  signal type_cast_327_inst_ack_0 : boolean;
  signal type_cast_327_inst_req_1 : boolean;
  signal type_cast_327_inst_ack_1 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal type_cast_328_inst_req_1 : boolean;
  signal type_cast_328_inst_ack_1 : boolean;
  signal addr_of_333_final_reg_req_0 : boolean;
  signal addr_of_333_final_reg_ack_0 : boolean;
  signal addr_of_333_final_reg_req_1 : boolean;
  signal addr_of_333_final_reg_ack_1 : boolean;
  signal ptr_deref_336_store_0_req_0 : boolean;
  signal ptr_deref_336_store_0_ack_0 : boolean;
  signal ptr_deref_336_store_0_req_1 : boolean;
  signal ptr_deref_336_store_0_ack_1 : boolean;
  signal ptr_deref_343_load_0_req_0 : boolean;
  signal ptr_deref_343_load_0_ack_0 : boolean;
  signal ptr_deref_343_load_0_req_1 : boolean;
  signal ptr_deref_343_load_0_ack_1 : boolean;
  signal ADD_u16_u16_349_inst_req_0 : boolean;
  signal ADD_u16_u16_349_inst_ack_0 : boolean;
  signal ADD_u16_u16_349_inst_req_1 : boolean;
  signal ADD_u16_u16_349_inst_ack_1 : boolean;
  signal ptr_deref_352_store_0_req_0 : boolean;
  signal ptr_deref_352_store_0_ack_0 : boolean;
  signal ptr_deref_352_store_0_req_1 : boolean;
  signal ptr_deref_352_store_0_ack_1 : boolean;
  signal RPIPE_rate_in_358_inst_req_0 : boolean;
  signal RPIPE_rate_in_358_inst_ack_0 : boolean;
  signal RPIPE_rate_in_358_inst_req_1 : boolean;
  signal RPIPE_rate_in_358_inst_ack_1 : boolean;
  signal ptr_deref_361_store_0_req_0 : boolean;
  signal ptr_deref_361_store_0_ack_0 : boolean;
  signal ptr_deref_361_store_0_req_1 : boolean;
  signal ptr_deref_361_store_0_ack_1 : boolean;
  signal ptr_deref_366_load_0_req_0 : boolean;
  signal ptr_deref_366_load_0_ack_0 : boolean;
  signal ptr_deref_366_load_0_req_1 : boolean;
  signal ptr_deref_366_load_0_ack_1 : boolean;
  signal STORE_rate_368_store_0_req_0 : boolean;
  signal STORE_rate_368_store_0_ack_0 : boolean;
  signal STORE_rate_368_store_0_req_1 : boolean;
  signal STORE_rate_368_store_0_ack_1 : boolean;
  signal memory_space_10_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_10_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_10_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_11_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_11_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_11_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_12_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_12_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_12_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_12_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_12_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_12_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_13_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_13_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_13_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_13_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_13_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_14_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_14_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_14_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_14_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_14_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_14_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_14_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initInputs_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initInputs_CP_117_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initInputs_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initInputs_CP_117_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initInputs_CP_117_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initInputs_CP_117_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initInputs_CP_117: Block -- control-path 
    signal initInputs_CP_117_elements: BooleanArray(237 downto 0);
    -- 
  begin -- 
    initInputs_CP_117_elements(0) <= initInputs_CP_117_start;
    initInputs_CP_117_symbol <= initInputs_CP_117_elements(237);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_43/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	27 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_43/branch_block_stmt_43__entry__
      -- CP-element group 1: 	 branch_block_stmt_43/assign_stmt_53_to_assign_stmt_73__entry__
      -- 
    initInputs_CP_117_elements(1) <= initInputs_CP_117_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	27 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_53_to_assign_stmt_73__exit__
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_76__entry__
      -- 
    initInputs_CP_117_elements(2) <= initInputs_CP_117_elements(27);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	30 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	31 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_76__exit__
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87__entry__
      -- 
    initInputs_CP_117_elements(3) <= initInputs_CP_117_elements(30);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	41 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	42 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87__exit__
      -- CP-element group 4: 	 branch_block_stmt_43/assign_stmt_90__entry__
      -- 
    initInputs_CP_117_elements(4) <= initInputs_CP_117_elements(41);
    -- CP-element group 5:  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	44 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	45 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_43/assign_stmt_90__exit__
      -- CP-element group 5: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106__entry__
      -- 
    initInputs_CP_117_elements(5) <= initInputs_CP_117_elements(44);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	57 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	208 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106__exit__
      -- CP-element group 6: 	 branch_block_stmt_43/bb_0_bb_1
      -- 
    initInputs_CP_117_elements(6) <= initInputs_CP_117_elements(57);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	211 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	58 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_43/merge_stmt_108__exit__
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127__entry__
      -- 
    initInputs_CP_117_elements(7) <= initInputs_CP_117_elements(211);
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	64 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	65 
    -- CP-element group 8: 	66 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127__exit__
      -- CP-element group 8: 	 branch_block_stmt_43/if_stmt_128__entry__
      -- 
    initInputs_CP_117_elements(8) <= initInputs_CP_117_elements(64);
    -- CP-element group 9:  merge  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	214 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	74 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_43/merge_stmt_134__exit__
      -- CP-element group 9: 	 branch_block_stmt_43/assign_stmt_137__entry__
      -- 
    initInputs_CP_117_elements(9) <= initInputs_CP_117_elements(214);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	76 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	77 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_137__exit__
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163__entry__
      -- 
    initInputs_CP_117_elements(10) <= initInputs_CP_117_elements(76);
    -- CP-element group 11:  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	93 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	215 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163__exit__
      -- CP-element group 11: 	 branch_block_stmt_43/bb_2_bb_3
      -- 
    initInputs_CP_117_elements(11) <= initInputs_CP_117_elements(93);
    -- CP-element group 12:  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	217 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	94 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_43/merge_stmt_165__exit__
      -- CP-element group 12: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179__entry__
      -- 
    initInputs_CP_117_elements(12) <= initInputs_CP_117_elements(217);
    -- CP-element group 13:  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	101 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	209 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179__exit__
      -- CP-element group 13: 	 branch_block_stmt_43/bb_3_bb_1
      -- 
    initInputs_CP_117_elements(13) <= initInputs_CP_117_elements(101);
    -- CP-element group 14:  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	220 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	103 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_43/merge_stmt_181__exit__
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266__entry__
      -- 
    initInputs_CP_117_elements(14) <= initInputs_CP_117_elements(220);
    -- CP-element group 15:  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	137 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	221 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266__exit__
      -- CP-element group 15: 	 branch_block_stmt_43/bb_4_bb_5
      -- 
    initInputs_CP_117_elements(15) <= initInputs_CP_117_elements(137);
    -- CP-element group 16:  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	224 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	138 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_43/merge_stmt_268__exit__
      -- CP-element group 16: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291__entry__
      -- 
    initInputs_CP_117_elements(16) <= initInputs_CP_117_elements(224);
    -- CP-element group 17:  branch  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	149 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	150 
    -- CP-element group 17: 	151 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291__exit__
      -- CP-element group 17: 	 branch_block_stmt_43/if_stmt_292__entry__
      -- 
    initInputs_CP_117_elements(17) <= initInputs_CP_117_elements(149);
    -- CP-element group 18:  merge  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	227 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	159 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_43/merge_stmt_298__exit__
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_301__entry__
      -- 
    initInputs_CP_117_elements(18) <= initInputs_CP_117_elements(227);
    -- CP-element group 19:  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	161 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	162 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_301__exit__
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338__entry__
      -- 
    initInputs_CP_117_elements(19) <= initInputs_CP_117_elements(161);
    -- CP-element group 20:  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	184 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	228 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338__exit__
      -- CP-element group 20: 	 branch_block_stmt_43/bb_6_bb_7
      -- 
    initInputs_CP_117_elements(20) <= initInputs_CP_117_elements(184);
    -- CP-element group 21:  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	230 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	185 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_43/merge_stmt_340__exit__
      -- CP-element group 21: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354__entry__
      -- 
    initInputs_CP_117_elements(21) <= initInputs_CP_117_elements(230);
    -- CP-element group 22:  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	192 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	222 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354__exit__
      -- CP-element group 22: 	 branch_block_stmt_43/bb_7_bb_5
      -- 
    initInputs_CP_117_elements(22) <= initInputs_CP_117_elements(192);
    -- CP-element group 23:  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	233 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	194 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_43/merge_stmt_356__exit__
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_359__entry__
      -- 
    initInputs_CP_117_elements(23) <= initInputs_CP_117_elements(233);
    -- CP-element group 24:  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	196 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	197 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_43/assign_stmt_359__exit__
      -- CP-element group 24: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370__entry__
      -- 
    initInputs_CP_117_elements(24) <= initInputs_CP_117_elements(196);
    -- CP-element group 25:  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	207 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	234 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370__exit__
      -- CP-element group 25: 	 branch_block_stmt_43/return__
      -- 
    initInputs_CP_117_elements(25) <= initInputs_CP_117_elements(207);
    -- CP-element group 26:  place  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	236 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	237 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_43/branch_block_stmt_43__exit__
      -- CP-element group 26: 	 branch_block_stmt_43/merge_stmt_372__exit__
      -- 
    initInputs_CP_117_elements(26) <= initInputs_CP_117_elements(236);
    -- CP-element group 27:  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	2 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_53_to_assign_stmt_73/$entry
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_53_to_assign_stmt_73/$exit
      -- 
    initInputs_CP_117_elements(27) <= initInputs_CP_117_elements(1);
    -- CP-element group 28:  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_76/$entry
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Sample/rr
      -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(28), ack => RPIPE_maxNitr_in_75_inst_req_0); -- 
    initInputs_CP_117_elements(28) <= initInputs_CP_117_elements(2);
    -- CP-element group 29:  transition  input  output  no-bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_update_start_
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Update/cr
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxNitr_in_75_inst_ack_0, ack => initInputs_CP_117_elements(29)); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(29), ack => RPIPE_maxNitr_in_75_inst_req_1); -- 
    -- CP-element group 30:  transition  input  no-bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	3 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_76/$exit
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_76/RPIPE_maxNitr_in_75_Update/ca
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxNitr_in_75_inst_ack_1, ack => initInputs_CP_117_elements(30)); -- 
    -- CP-element group 31:  fork  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	3 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	39 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	34 
    -- CP-element group 31: 	37 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (59) 
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/word_0/cr
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_update_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_address_resized
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_addr_resize/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_addr_resize/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_addr_resize/base_resize_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_addr_resize/base_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_word_addrgen/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_word_addrgen/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_word_addrgen/root_register_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_word_addrgen/root_register_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/ptr_deref_78_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/ptr_deref_78_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/ptr_deref_78_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/ptr_deref_78_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/word_0/cr
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_update_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_address_resized
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_addr_resize/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_addr_resize/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_addr_resize/base_resize_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_addr_resize/base_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_word_addrgen/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_word_addrgen/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_word_addrgen/root_register_req
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_word_addrgen/root_register_ack
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_update_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/word_0/cr
      -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(31), ack => ptr_deref_83_load_0_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(31), ack => ptr_deref_78_store_0_req_1); -- 
    rr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(31), ack => ptr_deref_78_store_0_req_0); -- 
    cr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(31), ack => STORE_maxNitr_85_store_0_req_1); -- 
    initInputs_CP_117_elements(31) <= initInputs_CP_117_elements(3);
    -- CP-element group 32:  transition  input  no-bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	40 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Sample/word_access_start/word_0/ra
      -- 
    ra_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_78_store_0_ack_0, ack => initInputs_CP_117_elements(32)); -- 
    -- CP-element group 33:  transition  input  no-bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	41 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_Update/word_access_complete/word_0/ca
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_78_store_0_ack_1, ack => initInputs_CP_117_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/word_0/rr
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/$entry
      -- 
    rr_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(34), ack => ptr_deref_83_load_0_req_0); -- 
    initInputs_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(40) & initInputs_CP_117_elements(31);
      gj_initInputs_cp_element_group_34 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  no-bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/word_0/ra
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Sample/word_access_start/$exit
      -- 
    ra_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_83_load_0_ack_0, ack => initInputs_CP_117_elements(35)); -- 
    -- CP-element group 36:  transition  input  no-bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/word_access_complete/word_0/ca
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/ptr_deref_83_Merge/$entry
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/ptr_deref_83_Merge/$exit
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/ptr_deref_83_Merge/merge_req
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_Update/ptr_deref_83_Merge/merge_ack
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_83_update_completed_
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_83_load_0_ack_1, ack => initInputs_CP_117_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	31 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/STORE_maxNitr_85_Split/$entry
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/STORE_maxNitr_85_Split/$exit
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/STORE_maxNitr_85_Split/split_req
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/STORE_maxNitr_85_Split/split_ack
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/word_0/rr
      -- 
    rr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(37), ack => STORE_maxNitr_85_store_0_req_0); -- 
    initInputs_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(31) & initInputs_CP_117_elements(36);
      gj_initInputs_cp_element_group_37 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  no-bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Sample/word_access_start/word_0/ra
      -- 
    ra_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_maxNitr_85_store_0_ack_0, ack => initInputs_CP_117_elements(38)); -- 
    -- CP-element group 39:  transition  input  no-bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	31 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/STORE_maxNitr_85_Update/word_access_complete/word_0/ca
      -- 
    ca_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_maxNitr_85_store_0_ack_1, ack => initInputs_CP_117_elements(39)); -- 
    -- CP-element group 40:  transition  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	32 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	34 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/ptr_deref_78_ptr_deref_83_delay
      -- 
    -- Element group initInputs_CP_117_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(32), ack => initInputs_CP_117_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	33 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	4 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_43/assign_stmt_80_to_assign_stmt_87/$exit
      -- 
    initInputs_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(39) & initInputs_CP_117_elements(33);
      gj_initInputs_cp_element_group_41 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	4 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_90/$entry
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Sample/rr
      -- 
    rr_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(42), ack => RPIPE_ebbyNo_in_89_inst_req_0); -- 
    initInputs_CP_117_elements(42) <= initInputs_CP_117_elements(4);
    -- CP-element group 43:  transition  input  output  no-bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_update_start_
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Update/cr
      -- 
    ra_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ebbyNo_in_89_inst_ack_0, ack => initInputs_CP_117_elements(43)); -- 
    cr_351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(43), ack => RPIPE_ebbyNo_in_89_inst_req_1); -- 
    -- CP-element group 44:  transition  input  no-bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	5 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_90/$exit
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_90/RPIPE_ebbyNo_in_89_Update/ca
      -- 
    ca_352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ebbyNo_in_89_inst_ack_1, ack => initInputs_CP_117_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	5 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	48 
    -- CP-element group 45: 	50 
    -- CP-element group 45: 	51 
    -- CP-element group 45: 	53 
    -- CP-element group 45: 	54 
    -- CP-element group 45: 	55 
    -- CP-element group 45:  members (89) 
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_update_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_word_addrgen/root_register_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/ptr_deref_92_Split/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/ptr_deref_92_Split/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/ptr_deref_92_Split/split_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/ptr_deref_92_Split/split_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/word_0/rr
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/word_0/cr
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_update_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_word_addrgen/root_register_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/word_0/cr
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_update_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/word_0/cr
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_update_start_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_word_addrgen/root_register_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/ptr_deref_103_Split/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/ptr_deref_103_Split/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/ptr_deref_103_Split/split_req
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/ptr_deref_103_Split/split_ack
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/word_0/rr
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/word_0/cr
      -- 
    cr_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => ptr_deref_97_load_0_req_1); -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => STORE_ebbyNo_99_store_0_req_1); -- 
    cr_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => ptr_deref_103_store_0_req_1); -- 
    rr_526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => ptr_deref_103_store_0_req_0); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => ptr_deref_92_store_0_req_1); -- 
    rr_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(45), ack => ptr_deref_92_store_0_req_0); -- 
    initInputs_CP_117_elements(45) <= initInputs_CP_117_elements(5);
    -- CP-element group 46:  transition  input  no-bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	56 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Sample/word_access_start/word_0/ra
      -- 
    ra_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_92_store_0_ack_0, ack => initInputs_CP_117_elements(46)); -- 
    -- CP-element group 47:  transition  input  no-bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	57 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_Update/word_access_complete/word_0/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_92_store_0_ack_1, ack => initInputs_CP_117_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	56 
    -- CP-element group 48: 	45 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/word_0/rr
      -- 
    rr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(48), ack => ptr_deref_97_load_0_req_0); -- 
    initInputs_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(56) & initInputs_CP_117_elements(45);
      gj_initInputs_cp_element_group_48 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  no-bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Sample/word_access_start/word_0/ra
      -- 
    ra_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_97_load_0_ack_0, ack => initInputs_CP_117_elements(49)); -- 
    -- CP-element group 50:  transition  input  no-bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/word_access_complete/word_0/ca
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/ptr_deref_97_Merge/$entry
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/ptr_deref_97_Merge/$exit
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/ptr_deref_97_Merge/merge_req
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_97_Update/ptr_deref_97_Merge/merge_ack
      -- 
    ca_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_97_load_0_ack_1, ack => initInputs_CP_117_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: 	45 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/STORE_ebbyNo_99_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/STORE_ebbyNo_99_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/STORE_ebbyNo_99_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/STORE_ebbyNo_99_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/word_0/rr
      -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(51), ack => STORE_ebbyNo_99_store_0_req_0); -- 
    initInputs_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(50) & initInputs_CP_117_elements(45);
      gj_initInputs_cp_element_group_51 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  no-bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Sample/word_access_start/word_0/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ebbyNo_99_store_0_ack_0, ack => initInputs_CP_117_elements(52)); -- 
    -- CP-element group 53:  transition  input  no-bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	45 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/STORE_ebbyNo_99_Update/word_access_complete/word_0/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ebbyNo_99_store_0_ack_1, ack => initInputs_CP_117_elements(53)); -- 
    -- CP-element group 54:  transition  input  no-bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	45 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Sample/word_access_start/word_0/ra
      -- 
    ra_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_103_store_0_ack_0, ack => initInputs_CP_117_elements(54)); -- 
    -- CP-element group 55:  transition  input  no-bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	45 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_103_Update/word_access_complete/word_0/ca
      -- 
    ca_538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_103_store_0_ack_1, ack => initInputs_CP_117_elements(55)); -- 
    -- CP-element group 56:  transition  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	46 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	48 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/ptr_deref_92_ptr_deref_97_delay
      -- 
    -- Element group initInputs_CP_117_elements(56) is a control-delay.
    cp_element_56_delay: control_delay_element  generic map(name => " 56_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(46), ack => initInputs_CP_117_elements(56), clk => clk, reset =>reset);
    -- CP-element group 57:  join  transition  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	47 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	6 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_43/assign_stmt_94_to_assign_stmt_106/$exit
      -- 
    initInputs_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(47) & initInputs_CP_117_elements(53) & initInputs_CP_117_elements(55);
      gj_initInputs_cp_element_group_57 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  fork  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	7 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (33) 
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_update_start_
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/word_0/rr
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_update_start_
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_update_start_
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Update/cr
      -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(58), ack => ptr_deref_111_load_0_req_1); -- 
    rr_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(58), ack => ptr_deref_111_load_0_req_0); -- 
    cr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(58), ack => type_cast_116_inst_req_1); -- 
    cr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(58), ack => SLT_i32_u1_125_inst_req_1); -- 
    initInputs_CP_117_elements(58) <= initInputs_CP_117_elements(7);
    -- CP-element group 59:  transition  input  no-bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Sample/word_access_start/word_0/ra
      -- 
    ra_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_111_load_0_ack_0, ack => initInputs_CP_117_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  no-bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/ptr_deref_111_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/ptr_deref_111_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/ptr_deref_111_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/ptr_deref_111_Update/ptr_deref_111_Merge/merge_ack
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Sample/rr
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_111_load_0_ack_1, ack => initInputs_CP_117_elements(60)); -- 
    rr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(60), ack => type_cast_116_inst_req_0); -- 
    -- CP-element group 61:  transition  input  no-bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Sample/ra
      -- 
    ra_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_116_inst_ack_0, ack => initInputs_CP_117_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  no-bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/type_cast_116_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Sample/rr
      -- 
    ca_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_116_inst_ack_1, ack => initInputs_CP_117_elements(62)); -- 
    rr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(62), ack => SLT_i32_u1_125_inst_req_0); -- 
    -- CP-element group 63:  transition  input  no-bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Sample/ra
      -- 
    ra_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_125_inst_ack_0, ack => initInputs_CP_117_elements(63)); -- 
    -- CP-element group 64:  transition  input  no-bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	8 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/$exit
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_112_to_assign_stmt_127/SLT_i32_u1_125_Update/ca
      -- 
    ca_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_125_inst_ack_1, ack => initInputs_CP_117_elements(64)); -- 
    -- CP-element group 65:  transition  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	8 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_43/if_stmt_128_dead_link/$entry
      -- 
    initInputs_CP_117_elements(65) <= initInputs_CP_117_elements(8);
    -- CP-element group 66:  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	8 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_43/if_stmt_128_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_43/if_stmt_128_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_43/if_stmt_128_eval_test/branch_req
      -- 
    branch_req_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(66), ack => if_stmt_128_branch_req_0); -- 
    initInputs_CP_117_elements(66) <= initInputs_CP_117_elements(8);
    -- CP-element group 67:  branch  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_43/R_iNsTr_14_129_place
      -- 
    initInputs_CP_117_elements(67) <= initInputs_CP_117_elements(66);
    -- CP-element group 68:  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_43/if_stmt_128_if_link/$entry
      -- 
    initInputs_CP_117_elements(68) <= initInputs_CP_117_elements(67);
    -- CP-element group 69:  transition  input  no-bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	72 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_43/if_stmt_128_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_43/if_stmt_128_if_link/if_choice_transition
      -- 
    if_choice_transition_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_128_branch_ack_1, ack => initInputs_CP_117_elements(69)); -- 
    -- CP-element group 70:  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_43/if_stmt_128_else_link/$entry
      -- 
    initInputs_CP_117_elements(70) <= initInputs_CP_117_elements(67);
    -- CP-element group 71:  transition  input  no-bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_43/if_stmt_128_else_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_43/if_stmt_128_else_link/else_choice_transition
      -- 
    else_choice_transition_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_128_branch_ack_0, ack => initInputs_CP_117_elements(71)); -- 
    -- CP-element group 72:  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	69 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	212 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_43/bb_1_bb_2
      -- 
    initInputs_CP_117_elements(72) <= initInputs_CP_117_elements(69);
    -- CP-element group 73:  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	218 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_43/bb_1_bb_4
      -- 
    initInputs_CP_117_elements(73) <= initInputs_CP_117_elements(71);
    -- CP-element group 74:  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	9 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_137/$entry
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Sample/rr
      -- 
    rr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(74), ack => RPIPE_matrix_in_136_inst_req_0); -- 
    initInputs_CP_117_elements(74) <= initInputs_CP_117_elements(9);
    -- CP-element group 75:  transition  input  output  no-bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (6) 
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_update_start_
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Update/cr
      -- 
    ra_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_136_inst_ack_0, ack => initInputs_CP_117_elements(75)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(75), ack => RPIPE_matrix_in_136_inst_req_1); -- 
    -- CP-element group 76:  transition  input  no-bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	10 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_137/$exit
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_137/RPIPE_matrix_in_136_Update/ca
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_136_inst_ack_1, ack => initInputs_CP_117_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	10 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	80 
    -- CP-element group 77: 	82 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	86 
    -- CP-element group 77: 	88 
    -- CP-element group 77: 	91 
    -- CP-element group 77:  members (89) 
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/ptr_deref_139_Split/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/ptr_deref_139_Split/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/ptr_deref_139_Split/split_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/ptr_deref_139_Split/split_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_complete/req
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_update_start_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/word_0/cr
      -- 
    cr_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_139_store_0_req_1); -- 
    rr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_139_store_0_req_0); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_144_load_0_req_1); -- 
    cr_803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_148_load_0_req_1); -- 
    rr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_148_load_0_req_0); -- 
    cr_822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => type_cast_153_inst_req_1); -- 
    req_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => addr_of_158_final_reg_req_1); -- 
    cr_911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(77), ack => ptr_deref_161_store_0_req_1); -- 
    initInputs_CP_117_elements(77) <= initInputs_CP_117_elements(10);
    -- CP-element group 78:  transition  input  no-bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	92 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/$exit
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Sample/word_access_start/word_0/ra
      -- 
    ra_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_store_0_ack_0, ack => initInputs_CP_117_elements(78)); -- 
    -- CP-element group 79:  transition  input  no-bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	93 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_Update/word_access_complete/word_0/ca
      -- 
    ca_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_store_0_ack_1, ack => initInputs_CP_117_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: 	92 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/word_0/rr
      -- 
    rr_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(80), ack => ptr_deref_144_load_0_req_0); -- 
    initInputs_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(77) & initInputs_CP_117_elements(92);
      gj_initInputs_cp_element_group_80 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  no-bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Sample/word_access_start/word_0/ra
      -- 
    ra_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_144_load_0_ack_0, ack => initInputs_CP_117_elements(81)); -- 
    -- CP-element group 82:  transition  input  no-bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	77 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	89 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/word_access_complete/word_0/ca
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/ptr_deref_144_Merge/$entry
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/ptr_deref_144_Merge/$exit
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/ptr_deref_144_Merge/merge_req
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_144_Update/ptr_deref_144_Merge/merge_ack
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_144_load_0_ack_1, ack => initInputs_CP_117_elements(82)); -- 
    -- CP-element group 83:  transition  input  no-bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/$exit
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Sample/word_access_start/word_0/ra
      -- 
    ra_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_148_load_0_ack_0, ack => initInputs_CP_117_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  no-bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (12) 
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/word_access_complete/word_0/ca
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/ptr_deref_148_Merge/$entry
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/ptr_deref_148_Merge/$exit
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/ptr_deref_148_Merge/merge_req
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_148_Update/ptr_deref_148_Merge/merge_ack
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Sample/rr
      -- 
    ca_804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_148_load_0_ack_1, ack => initInputs_CP_117_elements(84)); -- 
    rr_817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(84), ack => type_cast_153_inst_req_0); -- 
    -- CP-element group 85:  transition  input  no-bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Sample/ra
      -- 
    ra_818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => initInputs_CP_117_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  no-bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	77 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (27) 
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/type_cast_153_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_root_address_calculated
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_offset_calculated
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_resized_0
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_scaled_0
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_computed_0
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_resize_0/$entry
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_resize_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_resize_0/index_resize_req
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_resize_0/index_resize_ack
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_scale_0/$entry
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_scale_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_scale_0/scale_rename_req
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_index_scale_0/scale_rename_ack
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_final_index_sum_regn/$entry
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_final_index_sum_regn/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_final_index_sum_regn/req
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_final_index_sum_regn/ack
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_base_plus_offset/$entry
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_base_plus_offset/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_base_plus_offset/sum_rename_req
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/array_obj_ref_157_base_plus_offset/sum_rename_ack
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_request/$entry
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_request/req
      -- 
    ca_823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => initInputs_CP_117_elements(86)); -- 
    req_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(86), ack => addr_of_158_final_reg_req_0); -- 
    -- CP-element group 87:  transition  input  no-bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_request/$exit
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_request/ack
      -- 
    ack_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_158_final_reg_ack_0, ack => initInputs_CP_117_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  no-bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	77 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (19) 
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_complete/$exit
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/addr_of_158_complete/ack
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_word_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_address_resized
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_addr_resize/$entry
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_addr_resize/$exit
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_addr_resize/base_resize_req
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_addr_resize/base_resize_ack
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_word_addrgen/$entry
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_word_addrgen/$exit
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_word_addrgen/root_register_req
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_word_addrgen/root_register_ack
      -- 
    ack_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_158_final_reg_ack_1, ack => initInputs_CP_117_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	82 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/ptr_deref_161_Split/$entry
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/ptr_deref_161_Split/$exit
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/ptr_deref_161_Split/split_req
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/ptr_deref_161_Split/split_ack
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/word_0/rr
      -- 
    rr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(89), ack => ptr_deref_161_store_0_req_0); -- 
    initInputs_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(82) & initInputs_CP_117_elements(88);
      gj_initInputs_cp_element_group_89 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  no-bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/$exit
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Sample/word_access_start/word_0/ra
      -- 
    ra_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_161_store_0_ack_0, ack => initInputs_CP_117_elements(90)); -- 
    -- CP-element group 91:  transition  input  no-bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	77 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/$exit
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_161_Update/word_access_complete/word_0/ca
      -- 
    ca_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_161_store_0_ack_1, ack => initInputs_CP_117_elements(91)); -- 
    -- CP-element group 92:  transition  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	78 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	80 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/ptr_deref_139_ptr_deref_144_delay
      -- 
    -- Element group initInputs_CP_117_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(78), ack => initInputs_CP_117_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	79 
    -- CP-element group 93: 	87 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	11 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_43/assign_stmt_141_to_assign_stmt_163/$exit
      -- 
    initInputs_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(79) & initInputs_CP_117_elements(87) & initInputs_CP_117_elements(91);
      gj_initInputs_cp_element_group_93 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  fork  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	12 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	96 
    -- CP-element group 94: 	98 
    -- CP-element group 94: 	99 
    -- CP-element group 94: 	101 
    -- CP-element group 94:  members (51) 
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_update_start_
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_word_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_root_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_address_resized
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_addr_resize/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_addr_resize/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_addr_resize/base_resize_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_addr_resize/base_resize_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_plus_offset/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_plus_offset/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_plus_offset/sum_rename_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_base_plus_offset/sum_rename_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_word_addrgen/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_word_addrgen/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_word_addrgen/root_register_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_word_addrgen/root_register_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_update_start_
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_update_start_
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_word_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_root_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_address_resized
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_addr_resize/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_addr_resize/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_addr_resize/base_resize_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_addr_resize/base_resize_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_plus_offset/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_plus_offset/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_plus_offset/sum_rename_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_base_plus_offset/sum_rename_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_word_addrgen/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_word_addrgen/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_word_addrgen/root_register_req
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_word_addrgen/root_register_ack
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/word_0/cr
      -- 
    cr_960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(94), ack => ptr_deref_168_load_0_req_1); -- 
    rr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(94), ack => ptr_deref_168_load_0_req_0); -- 
    cr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(94), ack => ADD_u16_u16_174_inst_req_1); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(94), ack => ptr_deref_177_store_0_req_1); -- 
    initInputs_CP_117_elements(94) <= initInputs_CP_117_elements(12);
    -- CP-element group 95:  transition  input  no-bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	102 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Sample/word_access_start/word_0/ra
      -- 
    ra_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_168_load_0_ack_0, ack => initInputs_CP_117_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  no-bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (12) 
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/ptr_deref_168_Merge/$entry
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/ptr_deref_168_Merge/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/ptr_deref_168_Merge/merge_req
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_Update/ptr_deref_168_Merge/merge_ack
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Sample/rr
      -- 
    ca_961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_168_load_0_ack_1, ack => initInputs_CP_117_elements(96)); -- 
    rr_974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(96), ack => ADD_u16_u16_174_inst_req_0); -- 
    -- CP-element group 97:  transition  input  no-bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Sample/ra
      -- 
    ra_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_174_inst_ack_0, ack => initInputs_CP_117_elements(97)); -- 
    -- CP-element group 98:  transition  input  no-bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	94 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ADD_u16_u16_174_Update/ca
      -- 
    ca_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_174_inst_ack_1, ack => initInputs_CP_117_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  no-bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	94 
    -- CP-element group 99: 	98 
    -- CP-element group 99: 	102 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/ptr_deref_177_Split/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/ptr_deref_177_Split/$exit
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/ptr_deref_177_Split/split_req
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/ptr_deref_177_Split/split_ack
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/word_0/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/word_0/rr
      -- 
    rr_1018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(99), ack => ptr_deref_177_store_0_req_0); -- 
    initInputs_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(94) & initInputs_CP_117_elements(98) & initInputs_CP_117_elements(102);
      gj_initInputs_cp_element_group_99 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  transition  input  no-bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/$exit
      -- CP-element group 100: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Sample/word_access_start/word_0/ra
      -- 
    ra_1019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_177_store_0_ack_0, ack => initInputs_CP_117_elements(100)); -- 
    -- CP-element group 101:  transition  input  no-bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	94 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	13 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/$exit
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/$exit
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_177_Update/word_access_complete/word_0/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_177_store_0_ack_1, ack => initInputs_CP_117_elements(101)); -- 
    -- CP-element group 102:  transition  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	95 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	99 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_169_to_assign_stmt_179/ptr_deref_168_ptr_deref_177_delay
      -- 
    -- Element group initInputs_CP_117_elements(102) is a control-delay.
    cp_element_102_delay: control_delay_element  generic map(name => " 102_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(95), ack => initInputs_CP_117_elements(102), clk => clk, reset =>reset);
    -- CP-element group 103:  join  fork  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	14 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	105 
    -- CP-element group 103: 	106 
    -- CP-element group 103: 	108 
    -- CP-element group 103: 	109 
    -- CP-element group 103: 	110 
    -- CP-element group 103: 	111 
    -- CP-element group 103: 	113 
    -- CP-element group 103: 	114 
    -- CP-element group 103: 	115 
    -- CP-element group 103: 	116 
    -- CP-element group 103: 	118 
    -- CP-element group 103: 	119 
    -- CP-element group 103: 	120 
    -- CP-element group 103: 	122 
    -- CP-element group 103: 	123 
    -- CP-element group 103: 	124 
    -- CP-element group 103: 	126 
    -- CP-element group 103: 	129 
    -- CP-element group 103: 	131 
    -- CP-element group 103: 	132 
    -- CP-element group 103: 	134 
    -- CP-element group 103: 	135 
    -- CP-element group 103: 	136 
    -- CP-element group 103:  members (215) 
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/ptr_deref_263_Split/split_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/ptr_deref_263_Split/split_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/ptr_deref_263_Split/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/ptr_deref_263_Split/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_word_addrgen/root_register_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_word_addrgen/root_register_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/word_0/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/word_0/cr
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_update_start_
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_word_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_root_address_calculated
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_address_resized
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_addr_resize/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_addr_resize/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_addr_resize/base_resize_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_addr_resize/base_resize_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_plus_offset/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_plus_offset/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_plus_offset/sum_rename_req
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_base_plus_offset/sum_rename_ack
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_word_addrgen/$entry
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_word_addrgen/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_word_addrgen/root_register_req
      -- 
    cr_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_190_load_0_req_1); -- 
    rr_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_190_load_0_req_0); -- 
    cr_1116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => STORE_nrows_192_store_0_req_1); -- 
    cr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_203_load_0_req_1); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_203_load_0_req_0); -- 
    cr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => STORE_ncols_205_store_0_req_1); -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_216_load_0_req_1); -- 
    rr_1233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_216_load_0_req_0); -- 
    cr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => STORE_ncol_ind_218_store_0_req_1); -- 
    cr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_229_load_0_req_1); -- 
    rr_1316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_229_load_0_req_0); -- 
    cr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => type_cast_233_inst_req_1); -- 
    cr_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_243_load_0_req_1); -- 
    rr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_243_load_0_req_0); -- 
    cr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => type_cast_247_inst_req_1); -- 
    cr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ADD_u32_u32_252_inst_req_1); -- 
    cr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => type_cast_256_inst_req_1); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_259_store_0_req_1); -- 
    cr_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_263_store_0_req_1); -- 
    rr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(103), ack => ptr_deref_263_store_0_req_0); -- 
    initInputs_CP_117_elements(103) <= initInputs_CP_117_elements(14);
    -- CP-element group 104:  transition  input  no-bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/word_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Sample/word_access_start/word_0/ra
      -- 
    ra_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_load_0_ack_0, ack => initInputs_CP_117_elements(104)); -- 
    -- CP-element group 105:  transition  input  no-bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/$exit
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/word_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/word_access_complete/word_0/ca
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/ptr_deref_190_Merge/$entry
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/ptr_deref_190_Merge/$exit
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/ptr_deref_190_Merge/merge_req
      -- CP-element group 105: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_190_Update/ptr_deref_190_Merge/merge_ack
      -- 
    ca_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_load_0_ack_1, ack => initInputs_CP_117_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  no-bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/STORE_nrows_192_Split/$entry
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/STORE_nrows_192_Split/$exit
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/STORE_nrows_192_Split/split_req
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/STORE_nrows_192_Split/split_ack
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/$entry
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/word_0/rr
      -- 
    rr_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(106), ack => STORE_nrows_192_store_0_req_0); -- 
    initInputs_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(103) & initInputs_CP_117_elements(105);
      gj_initInputs_cp_element_group_106 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  no-bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Sample/word_access_start/word_0/ra
      -- 
    ra_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_nrows_192_store_0_ack_0, ack => initInputs_CP_117_elements(107)); -- 
    -- CP-element group 108:  transition  input  no-bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	103 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	137 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_nrows_192_Update/word_access_complete/word_0/ca
      -- 
    ca_1117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_nrows_192_store_0_ack_1, ack => initInputs_CP_117_elements(108)); -- 
    -- CP-element group 109:  transition  input  no-bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	103 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_sample_completed_
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_203_load_0_ack_0, ack => initInputs_CP_117_elements(109)); -- 
    -- CP-element group 110:  transition  input  no-bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/ptr_deref_203_Merge/merge_ack
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/ptr_deref_203_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/ptr_deref_203_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_Update/ptr_deref_203_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_203_update_completed_
      -- 
    ca_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_203_load_0_ack_1, ack => initInputs_CP_117_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  no-bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	103 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/word_0/rr
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/word_0/$entry
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/$entry
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/STORE_ncols_205_Split/split_ack
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/STORE_ncols_205_Split/split_req
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/STORE_ncols_205_Split/$exit
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/STORE_ncols_205_Split/$entry
      -- CP-element group 111: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/$entry
      -- 
    rr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(111), ack => STORE_ncols_205_store_0_req_0); -- 
    initInputs_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(103) & initInputs_CP_117_elements(110);
      gj_initInputs_cp_element_group_111 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  no-bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Sample/$exit
      -- 
    ra_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncols_205_store_0_ack_0, ack => initInputs_CP_117_elements(112)); -- 
    -- CP-element group 113:  transition  input  no-bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	103 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	137 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/word_access_complete/$exit
      -- CP-element group 113: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncols_205_update_completed_
      -- 
    ca_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncols_205_store_0_ack_1, ack => initInputs_CP_117_elements(113)); -- 
    -- CP-element group 114:  transition  input  no-bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	103 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/word_0/ra
      -- CP-element group 114: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/word_access_start/$exit
      -- CP-element group 114: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_sample_completed_
      -- 
    ra_1234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_216_load_0_ack_0, ack => initInputs_CP_117_elements(114)); -- 
    -- CP-element group 115:  transition  input  no-bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	103 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (9) 
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/ptr_deref_216_Merge/merge_ack
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/ptr_deref_216_Merge/merge_req
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/ptr_deref_216_Merge/$exit
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/ptr_deref_216_Merge/$entry
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/word_0/ca
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/word_0/$exit
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/word_access_complete/$exit
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_216_update_completed_
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_216_load_0_ack_1, ack => initInputs_CP_117_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  no-bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	103 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/STORE_ncol_ind_218_Split/split_ack
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/STORE_ncol_ind_218_Split/split_req
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/STORE_ncol_ind_218_Split/$exit
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/STORE_ncol_ind_218_Split/$entry
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_sample_start_
      -- 
    rr_1271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(116), ack => STORE_ncol_ind_218_store_0_req_0); -- 
    initInputs_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(103) & initInputs_CP_117_elements(115);
      gj_initInputs_cp_element_group_116 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  no-bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/word_0/ra
      -- CP-element group 117: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_sample_completed_
      -- 
    ra_1272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncol_ind_218_store_0_ack_0, ack => initInputs_CP_117_elements(117)); -- 
    -- CP-element group 118:  transition  input  no-bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	103 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	137 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/STORE_ncol_ind_218_update_completed_
      -- 
    ca_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncol_ind_218_store_0_ack_1, ack => initInputs_CP_117_elements(118)); -- 
    -- CP-element group 119:  transition  input  no-bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	103 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/word_0/ra
      -- CP-element group 119: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Sample/$exit
      -- 
    ra_1317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_229_load_0_ack_0, ack => initInputs_CP_117_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  no-bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	103 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (12) 
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/ptr_deref_229_Merge/merge_ack
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/ptr_deref_229_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/ptr_deref_229_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/ptr_deref_229_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_229_Update/$exit
      -- 
    ca_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_229_load_0_ack_1, ack => initInputs_CP_117_elements(120)); -- 
    rr_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(120), ack => type_cast_233_inst_req_0); -- 
    -- CP-element group 121:  transition  input  no-bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Sample/ra
      -- CP-element group 121: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_sample_completed_
      -- 
    ra_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_0, ack => initInputs_CP_117_elements(121)); -- 
    -- CP-element group 122:  transition  input  no-bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	103 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	127 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_233_update_completed_
      -- 
    ca_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_1, ack => initInputs_CP_117_elements(122)); -- 
    -- CP-element group 123:  transition  input  no-bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	103 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (5) 
      -- CP-element group 123: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/word_0/ra
      -- CP-element group 123: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/word_0/$exit
      -- CP-element group 123: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/word_access_start/$exit
      -- CP-element group 123: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Sample/$exit
      -- 
    ra_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_243_load_0_ack_0, ack => initInputs_CP_117_elements(123)); -- 
    -- CP-element group 124:  transition  input  output  no-bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	103 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (12) 
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/ptr_deref_243_Merge/merge_req
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/ptr_deref_243_Merge/$exit
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/ptr_deref_243_Merge/$entry
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/word_0/ca
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Sample/rr
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/ptr_deref_243_Merge/merge_ack
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/word_access_complete/$exit
      -- CP-element group 124: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_243_Update/$exit
      -- 
    ca_1392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_243_load_0_ack_1, ack => initInputs_CP_117_elements(124)); -- 
    rr_1405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(124), ack => type_cast_247_inst_req_0); -- 
    -- CP-element group 125:  transition  input  no-bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Sample/ra
      -- CP-element group 125: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_sample_completed_
      -- 
    ra_1406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_247_inst_ack_0, ack => initInputs_CP_117_elements(125)); -- 
    -- CP-element group 126:  transition  input  no-bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	103 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Update/ca
      -- CP-element group 126: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_247_update_completed_
      -- 
    ca_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_247_inst_ack_1, ack => initInputs_CP_117_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_sample_start_
      -- 
    rr_1419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(127), ack => ADD_u32_u32_252_inst_req_0); -- 
    initInputs_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(122) & initInputs_CP_117_elements(126);
      gj_initInputs_cp_element_group_127 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  no-bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_sample_completed_
      -- 
    ra_1420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_252_inst_ack_0, ack => initInputs_CP_117_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  no-bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	103 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ADD_u32_u32_252_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Sample/rr
      -- 
    ca_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_252_inst_ack_1, ack => initInputs_CP_117_elements(129)); -- 
    rr_1433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(129), ack => type_cast_256_inst_req_0); -- 
    -- CP-element group 130:  transition  input  no-bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Sample/ra
      -- 
    ra_1434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_0, ack => initInputs_CP_117_elements(130)); -- 
    -- CP-element group 131:  transition  input  no-bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	103 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/type_cast_256_Update/$exit
      -- 
    ca_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_1, ack => initInputs_CP_117_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  no-bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	103 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/word_0/rr
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/ptr_deref_259_Split/$entry
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/$entry
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/word_0/$entry
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/ptr_deref_259_Split/split_ack
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/ptr_deref_259_Split/split_req
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/ptr_deref_259_Split/$exit
      -- 
    rr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(132), ack => ptr_deref_259_store_0_req_0); -- 
    initInputs_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(103) & initInputs_CP_117_elements(131);
      gj_initInputs_cp_element_group_132 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  transition  input  no-bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/word_0/ra
      -- CP-element group 133: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/word_0/$exit
      -- CP-element group 133: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Sample/word_access_start/$exit
      -- 
    ra_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_259_store_0_ack_0, ack => initInputs_CP_117_elements(133)); -- 
    -- CP-element group 134:  transition  input  no-bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	103 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/word_0/ca
      -- CP-element group 134: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_259_Update/word_access_complete/word_0/$exit
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_259_store_0_ack_1, ack => initInputs_CP_117_elements(134)); -- 
    -- CP-element group 135:  transition  input  no-bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	103 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/word_0/ra
      -- CP-element group 135: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/word_access_start/$exit
      -- CP-element group 135: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Sample/$exit
      -- 
    ra_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_store_0_ack_0, ack => initInputs_CP_117_elements(135)); -- 
    -- CP-element group 136:  transition  input  no-bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	103 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/word_0/ca
      -- CP-element group 136: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/word_0/$exit
      -- CP-element group 136: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/word_access_complete/$exit
      -- CP-element group 136: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/ptr_deref_263_Update/$exit
      -- 
    ca_1539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_store_0_ack_1, ack => initInputs_CP_117_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	108 
    -- CP-element group 137: 	113 
    -- CP-element group 137: 	118 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	15 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_43/assign_stmt_187_to_assign_stmt_266/$exit
      -- 
    initInputs_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(108) & initInputs_CP_117_elements(113) & initInputs_CP_117_elements(118) & initInputs_CP_117_elements(134) & initInputs_CP_117_elements(136);
      gj_initInputs_cp_element_group_137 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	16 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	140 
    -- CP-element group 138: 	142 
    -- CP-element group 138: 	143 
    -- CP-element group 138: 	144 
    -- CP-element group 138: 	146 
    -- CP-element group 138: 	149 
    -- CP-element group 138:  members (62) 
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_addr_resize/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_addr_resize/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_addr_resize/base_resize_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_addr_resize/base_resize_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_root_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_address_resized
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_plus_offset/sum_rename_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/word_0/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/word_0/rr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_word_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_word_addrgen/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_word_addrgen/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_word_addrgen/root_register_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_word_addrgen/root_register_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_plus_offset/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_plus_offset/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_base_plus_offset/sum_rename_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/word_0/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_update_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/word_0/cr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_update_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Update/cr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_update_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_word_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_root_address_calculated
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_address_resized
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_addr_resize/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_addr_resize/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_addr_resize/base_resize_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_addr_resize/base_resize_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_plus_offset/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_plus_offset/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_plus_offset/sum_rename_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_base_plus_offset/sum_rename_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_word_addrgen/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_word_addrgen/$exit
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_word_addrgen/root_register_req
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_word_addrgen/root_register_ack
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/word_0/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/word_0/rr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/word_0/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/word_0/cr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_update_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Update/cr
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_update_start_
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Update/cr
      -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => ptr_deref_271_load_0_req_1); -- 
    rr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => ptr_deref_271_load_0_req_0); -- 
    cr_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => type_cast_275_inst_req_1); -- 
    cr_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => ptr_deref_279_load_0_req_1); -- 
    rr_1639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => ptr_deref_279_load_0_req_0); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => type_cast_283_inst_req_1); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(138), ack => SLT_i32_u1_290_inst_req_1); -- 
    initInputs_CP_117_elements(138) <= initInputs_CP_117_elements(16);
    -- CP-element group 139:  transition  input  no-bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (5) 
      -- CP-element group 139: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/word_0/$exit
      -- CP-element group 139: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/word_0/ra
      -- CP-element group 139: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Sample/word_access_start/$exit
      -- 
    ra_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_271_load_0_ack_0, ack => initInputs_CP_117_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  no-bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (12) 
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/$exit
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/word_0/$exit
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/word_access_complete/word_0/ca
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/ptr_deref_271_Merge/$entry
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/ptr_deref_271_Merge/$exit
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/ptr_deref_271_Merge/merge_req
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_271_Update/ptr_deref_271_Merge/merge_ack
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Sample/rr
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_271_load_0_ack_1, ack => initInputs_CP_117_elements(140)); -- 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(140), ack => type_cast_275_inst_req_0); -- 
    -- CP-element group 141:  transition  input  no-bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Sample/ra
      -- 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_0, ack => initInputs_CP_117_elements(141)); -- 
    -- CP-element group 142:  transition  input  no-bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	138 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	147 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_275_Update/ca
      -- 
    ca_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_1, ack => initInputs_CP_117_elements(142)); -- 
    -- CP-element group 143:  transition  input  no-bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	138 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/$exit
      -- CP-element group 143: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Sample/word_access_start/word_0/ra
      -- 
    ra_1640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_279_load_0_ack_0, ack => initInputs_CP_117_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  no-bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	138 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (12) 
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/$exit
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/word_access_complete/word_0/ca
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/ptr_deref_279_Merge/$entry
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/ptr_deref_279_Merge/$exit
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/ptr_deref_279_Merge/merge_req
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/ptr_deref_279_Update/ptr_deref_279_Merge/merge_ack
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Sample/rr
      -- 
    ca_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_279_load_0_ack_1, ack => initInputs_CP_117_elements(144)); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(144), ack => type_cast_283_inst_req_0); -- 
    -- CP-element group 145:  transition  input  no-bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Sample/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_283_inst_ack_0, ack => initInputs_CP_117_elements(145)); -- 
    -- CP-element group 146:  transition  input  no-bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	138 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/type_cast_283_Update/ca
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_283_inst_ack_1, ack => initInputs_CP_117_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	142 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Sample/rr
      -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(147), ack => SLT_i32_u1_290_inst_req_0); -- 
    initInputs_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(142) & initInputs_CP_117_elements(146);
      gj_initInputs_cp_element_group_147 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  transition  input  no-bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_290_inst_ack_0, ack => initInputs_CP_117_elements(148)); -- 
    -- CP-element group 149:  transition  input  no-bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	138 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	17 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/$exit
      -- CP-element group 149: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_43/assign_stmt_272_to_assign_stmt_291/SLT_i32_u1_290_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_290_inst_ack_1, ack => initInputs_CP_117_elements(149)); -- 
    -- CP-element group 150:  transition  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	17 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_43/if_stmt_292_dead_link/$entry
      -- 
    initInputs_CP_117_elements(150) <= initInputs_CP_117_elements(17);
    -- CP-element group 151:  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	17 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_43/if_stmt_292_eval_test/$entry
      -- CP-element group 151: 	 branch_block_stmt_43/if_stmt_292_eval_test/$exit
      -- CP-element group 151: 	 branch_block_stmt_43/if_stmt_292_eval_test/branch_req
      -- 
    branch_req_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(151), ack => if_stmt_292_branch_req_0); -- 
    initInputs_CP_117_elements(151) <= initInputs_CP_117_elements(17);
    -- CP-element group 152:  branch  place  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (1) 
      -- CP-element group 152: 	 branch_block_stmt_43/R_iNsTr_53_293_place
      -- 
    initInputs_CP_117_elements(152) <= initInputs_CP_117_elements(151);
    -- CP-element group 153:  transition  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (1) 
      -- CP-element group 153: 	 branch_block_stmt_43/if_stmt_292_if_link/$entry
      -- 
    initInputs_CP_117_elements(153) <= initInputs_CP_117_elements(152);
    -- CP-element group 154:  transition  input  no-bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (2) 
      -- CP-element group 154: 	 branch_block_stmt_43/if_stmt_292_if_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_43/if_stmt_292_if_link/if_choice_transition
      -- 
    if_choice_transition_1697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_292_branch_ack_1, ack => initInputs_CP_117_elements(154)); -- 
    -- CP-element group 155:  transition  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	152 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_43/if_stmt_292_else_link/$entry
      -- 
    initInputs_CP_117_elements(155) <= initInputs_CP_117_elements(152);
    -- CP-element group 156:  transition  input  no-bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_43/if_stmt_292_else_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_43/if_stmt_292_else_link/else_choice_transition
      -- 
    else_choice_transition_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_292_branch_ack_0, ack => initInputs_CP_117_elements(156)); -- 
    -- CP-element group 157:  place  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	225 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_43/bb_5_bb_6
      -- 
    initInputs_CP_117_elements(157) <= initInputs_CP_117_elements(154);
    -- CP-element group 158:  place  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	231 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_43/bb_5_bb_8
      -- 
    initInputs_CP_117_elements(158) <= initInputs_CP_117_elements(156);
    -- CP-element group 159:  transition  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	18 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (4) 
      -- CP-element group 159: 	 branch_block_stmt_43/assign_stmt_301/$entry
      -- CP-element group 159: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Sample/rr
      -- 
    rr_1714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(159), ack => RPIPE_matrix_in_300_inst_req_0); -- 
    initInputs_CP_117_elements(159) <= initInputs_CP_117_elements(18);
    -- CP-element group 160:  transition  input  output  no-bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_update_start_
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Update/cr
      -- 
    ra_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_300_inst_ack_0, ack => initInputs_CP_117_elements(160)); -- 
    cr_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(160), ack => RPIPE_matrix_in_300_inst_req_1); -- 
    -- CP-element group 161:  transition  input  no-bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	19 
    -- CP-element group 161:  members (4) 
      -- CP-element group 161: 	 branch_block_stmt_43/assign_stmt_301/$exit
      -- CP-element group 161: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_43/assign_stmt_301/RPIPE_matrix_in_300_Update/ca
      -- 
    ca_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_300_inst_ack_1, ack => initInputs_CP_117_elements(161)); -- 
    -- CP-element group 162:  join  fork  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	19 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	165 
    -- CP-element group 162: 	167 
    -- CP-element group 162: 	168 
    -- CP-element group 162: 	169 
    -- CP-element group 162: 	171 
    -- CP-element group 162: 	173 
    -- CP-element group 162: 	175 
    -- CP-element group 162: 	177 
    -- CP-element group 162: 	179 
    -- CP-element group 162: 	182 
    -- CP-element group 162:  members (98) 
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_word_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_root_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_address_resized
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_addr_resize/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_addr_resize/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_addr_resize/base_resize_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_addr_resize/base_resize_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_plus_offset/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_plus_offset/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_plus_offset/sum_rename_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_base_plus_offset/sum_rename_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_word_addrgen/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_word_addrgen/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_word_addrgen/root_register_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_word_addrgen/root_register_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/ptr_deref_303_Split/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/ptr_deref_303_Split/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/ptr_deref_303_Split/split_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/ptr_deref_303_Split/split_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/word_0/rr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/word_0/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_word_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_root_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_address_resized
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_addr_resize/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_addr_resize/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_addr_resize/base_resize_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_addr_resize/base_resize_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_plus_offset/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_plus_offset/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_plus_offset/sum_rename_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_base_plus_offset/sum_rename_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_word_addrgen/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_word_addrgen/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_word_addrgen/root_register_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_word_addrgen/root_register_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/word_0/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_word_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_root_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_address_resized
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_addr_resize/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_addr_resize/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_addr_resize/base_resize_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_addr_resize/base_resize_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_plus_offset/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_plus_offset/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_plus_offset/sum_rename_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_base_plus_offset/sum_rename_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_word_addrgen/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_word_addrgen/$exit
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_word_addrgen/root_register_req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_word_addrgen/root_register_ack
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/word_0/rr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/word_0/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_complete/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_complete/req
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_update_start_
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/word_0/cr
      -- 
    cr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_303_store_0_req_1); -- 
    rr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_303_store_0_req_0); -- 
    cr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_308_load_0_req_1); -- 
    cr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_312_load_0_req_1); -- 
    rr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_312_load_0_req_0); -- 
    cr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => type_cast_316_inst_req_1); -- 
    cr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ADD_u32_u32_322_inst_req_1); -- 
    cr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => type_cast_328_inst_req_1); -- 
    cr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => type_cast_327_inst_req_1); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => addr_of_333_final_reg_req_1); -- 
    cr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(162), ack => ptr_deref_336_store_0_req_1); -- 
    initInputs_CP_117_elements(162) <= initInputs_CP_117_elements(19);
    -- CP-element group 163:  transition  input  no-bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	183 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/$exit
      -- CP-element group 163: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Sample/word_access_start/word_0/ra
      -- 
    ra_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_0, ack => initInputs_CP_117_elements(163)); -- 
    -- CP-element group 164:  transition  input  no-bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	184 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/$exit
      -- CP-element group 164: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_Update/word_access_complete/word_0/ca
      -- 
    ca_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_1, ack => initInputs_CP_117_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: 	183 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/$entry
      -- CP-element group 165: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/word_0/$entry
      -- CP-element group 165: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/word_0/rr
      -- 
    rr_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(165), ack => ptr_deref_308_load_0_req_0); -- 
    initInputs_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(162) & initInputs_CP_117_elements(183);
      gj_initInputs_cp_element_group_165 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  no-bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/$exit
      -- CP-element group 166: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/word_0/$exit
      -- CP-element group 166: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Sample/word_access_start/word_0/ra
      -- 
    ra_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_308_load_0_ack_0, ack => initInputs_CP_117_elements(166)); -- 
    -- CP-element group 167:  transition  input  no-bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	162 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	180 
    -- CP-element group 167:  members (9) 
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/$exit
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/word_0/$exit
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/word_access_complete/word_0/ca
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/ptr_deref_308_Merge/$entry
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/ptr_deref_308_Merge/$exit
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/ptr_deref_308_Merge/merge_req
      -- CP-element group 167: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_308_Update/ptr_deref_308_Merge/merge_ack
      -- 
    ca_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_308_load_0_ack_1, ack => initInputs_CP_117_elements(167)); -- 
    -- CP-element group 168:  transition  input  no-bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	162 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/$exit
      -- CP-element group 168: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/word_0/$exit
      -- CP-element group 168: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Sample/word_access_start/word_0/ra
      -- 
    ra_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_312_load_0_ack_0, ack => initInputs_CP_117_elements(168)); -- 
    -- CP-element group 169:  transition  input  output  no-bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	162 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (12) 
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/$exit
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/word_0/$exit
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/word_access_complete/word_0/ca
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/ptr_deref_312_Merge/$entry
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/ptr_deref_312_Merge/$exit
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/ptr_deref_312_Merge/merge_req
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_312_Update/ptr_deref_312_Merge/merge_ack
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Sample/rr
      -- 
    ca_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_312_load_0_ack_1, ack => initInputs_CP_117_elements(169)); -- 
    rr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(169), ack => type_cast_316_inst_req_0); -- 
    -- CP-element group 170:  transition  input  no-bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Sample/ra
      -- 
    ra_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_0, ack => initInputs_CP_117_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  no-bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	162 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_316_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Sample/rr
      -- 
    ca_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_316_inst_ack_1, ack => initInputs_CP_117_elements(171)); -- 
    rr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(171), ack => ADD_u32_u32_322_inst_req_0); -- 
    -- CP-element group 172:  transition  input  no-bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Sample/ra
      -- 
    ra_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_322_inst_ack_0, ack => initInputs_CP_117_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  no-bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	162 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ADD_u32_u32_322_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Sample/rr
      -- 
    ca_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_322_inst_ack_1, ack => initInputs_CP_117_elements(173)); -- 
    rr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(173), ack => type_cast_327_inst_req_0); -- 
    -- CP-element group 174:  transition  input  no-bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Sample/ra
      -- 
    ra_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_0, ack => initInputs_CP_117_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  no-bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	162 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_327_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Sample/rr
      -- 
    ca_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_1, ack => initInputs_CP_117_elements(175)); -- 
    rr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(175), ack => type_cast_328_inst_req_0); -- 
    -- CP-element group 176:  transition  input  no-bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Sample/ra
      -- 
    ra_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_0, ack => initInputs_CP_117_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  no-bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	162 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (27) 
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/type_cast_328_Update/ca
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_root_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_offset_calculated
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_resized_0
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_scaled_0
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_computed_0
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_resize_0/$entry
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_resize_0/$exit
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_resize_0/index_resize_req
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_resize_0/index_resize_ack
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_scale_0/$entry
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_scale_0/$exit
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_scale_0/scale_rename_req
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_index_scale_0/scale_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_final_index_sum_regn/$entry
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_final_index_sum_regn/$exit
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_final_index_sum_regn/req
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_final_index_sum_regn/ack
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_base_plus_offset/$entry
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_base_plus_offset/$exit
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_base_plus_offset/sum_rename_req
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/array_obj_ref_332_base_plus_offset/sum_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_request/$entry
      -- CP-element group 177: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_request/req
      -- 
    ca_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_1, ack => initInputs_CP_117_elements(177)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(177), ack => addr_of_333_final_reg_req_0); -- 
    -- CP-element group 178:  transition  input  no-bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	184 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_request/$exit
      -- CP-element group 178: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_request/ack
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_333_final_reg_ack_0, ack => initInputs_CP_117_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  no-bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	162 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (19) 
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_complete/$exit
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/addr_of_333_complete/ack
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_address_calculated
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_word_address_calculated
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_root_address_calculated
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_address_resized
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_addr_resize/$entry
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_addr_resize/$exit
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_addr_resize/base_resize_req
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_addr_resize/base_resize_ack
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_plus_offset/$entry
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_plus_offset/$exit
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_plus_offset/sum_rename_req
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_base_plus_offset/sum_rename_ack
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_word_addrgen/$entry
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_word_addrgen/$exit
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_word_addrgen/root_register_req
      -- CP-element group 179: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_word_addrgen/root_register_ack
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_333_final_reg_ack_1, ack => initInputs_CP_117_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	167 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/ptr_deref_336_Split/$entry
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/ptr_deref_336_Split/$exit
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/ptr_deref_336_Split/split_req
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/ptr_deref_336_Split/split_ack
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/$entry
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/word_0/$entry
      -- CP-element group 180: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/word_0/rr
      -- 
    rr_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(180), ack => ptr_deref_336_store_0_req_0); -- 
    initInputs_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(167) & initInputs_CP_117_elements(179);
      gj_initInputs_cp_element_group_180 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  transition  input  no-bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/$exit
      -- CP-element group 181: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Sample/word_access_start/word_0/ra
      -- 
    ra_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_336_store_0_ack_0, ack => initInputs_CP_117_elements(181)); -- 
    -- CP-element group 182:  transition  input  no-bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	162 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/$exit
      -- CP-element group 182: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/word_0/$exit
      -- CP-element group 182: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_336_Update/word_access_complete/word_0/ca
      -- 
    ca_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_336_store_0_ack_1, ack => initInputs_CP_117_elements(182)); -- 
    -- CP-element group 183:  transition  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	163 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	165 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/ptr_deref_303_ptr_deref_308_delay
      -- 
    -- Element group initInputs_CP_117_elements(183) is a control-delay.
    cp_element_183_delay: control_delay_element  generic map(name => " 183_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(163), ack => initInputs_CP_117_elements(183), clk => clk, reset =>reset);
    -- CP-element group 184:  join  transition  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	164 
    -- CP-element group 184: 	178 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	20 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_43/assign_stmt_305_to_assign_stmt_338/$exit
      -- 
    initInputs_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(164) & initInputs_CP_117_elements(178) & initInputs_CP_117_elements(182);
      gj_initInputs_cp_element_group_184 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  fork  transition  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	21 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	189 
    -- CP-element group 185: 	190 
    -- CP-element group 185: 	192 
    -- CP-element group 185:  members (51) 
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_update_start_
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_word_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_root_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_address_resized
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_addr_resize/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_addr_resize/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_addr_resize/base_resize_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_addr_resize/base_resize_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_plus_offset/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_plus_offset/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_plus_offset/sum_rename_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_word_addrgen/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_word_addrgen/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_word_addrgen/root_register_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_word_addrgen/root_register_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/word_0/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/word_0/rr
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/word_0/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/word_0/cr
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_update_start_
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_update_start_
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_word_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_root_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_address_resized
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_addr_resize/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_addr_resize/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_addr_resize/base_resize_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_addr_resize/base_resize_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_plus_offset/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_plus_offset/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_plus_offset/sum_rename_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_base_plus_offset/sum_rename_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_word_addrgen/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_word_addrgen/$exit
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_word_addrgen/root_register_req
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_word_addrgen/root_register_ack
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/word_0/$entry
      -- CP-element group 185: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/word_0/cr
      -- 
    cr_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(185), ack => ptr_deref_343_load_0_req_1); -- 
    rr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(185), ack => ptr_deref_343_load_0_req_0); -- 
    cr_2085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(185), ack => ADD_u16_u16_349_inst_req_1); -- 
    cr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(185), ack => ptr_deref_352_store_0_req_1); -- 
    initInputs_CP_117_elements(185) <= initInputs_CP_117_elements(21);
    -- CP-element group 186:  transition  input  no-bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	193 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/$exit
      -- CP-element group 186: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Sample/word_access_start/word_0/ra
      -- 
    ra_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_load_0_ack_0, ack => initInputs_CP_117_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  no-bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (12) 
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/$exit
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/word_0/$exit
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/word_access_complete/word_0/ca
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/ptr_deref_343_Merge/$entry
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/ptr_deref_343_Merge/$exit
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/ptr_deref_343_Merge/merge_req
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_Update/ptr_deref_343_Merge/merge_ack
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Sample/rr
      -- 
    ca_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_load_0_ack_1, ack => initInputs_CP_117_elements(187)); -- 
    rr_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(187), ack => ADD_u16_u16_349_inst_req_0); -- 
    -- CP-element group 188:  transition  input  no-bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Sample/ra
      -- 
    ra_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_349_inst_ack_0, ack => initInputs_CP_117_elements(188)); -- 
    -- CP-element group 189:  transition  input  no-bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	185 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ADD_u16_u16_349_Update/ca
      -- 
    ca_2086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_349_inst_ack_1, ack => initInputs_CP_117_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  no-bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	185 
    -- CP-element group 190: 	189 
    -- CP-element group 190: 	193 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/ptr_deref_352_Split/$entry
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/ptr_deref_352_Split/$exit
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/ptr_deref_352_Split/split_req
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/ptr_deref_352_Split/split_ack
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/$entry
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/word_0/$entry
      -- CP-element group 190: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/word_0/rr
      -- 
    rr_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(190), ack => ptr_deref_352_store_0_req_0); -- 
    initInputs_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(185) & initInputs_CP_117_elements(189) & initInputs_CP_117_elements(193);
      gj_initInputs_cp_element_group_190 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  transition  input  no-bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/$exit
      -- CP-element group 191: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/word_0/$exit
      -- CP-element group 191: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Sample/word_access_start/word_0/ra
      -- 
    ra_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_352_store_0_ack_0, ack => initInputs_CP_117_elements(191)); -- 
    -- CP-element group 192:  transition  input  no-bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	185 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	22 
    -- CP-element group 192:  members (6) 
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/$exit
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/$exit
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/word_0/$exit
      -- CP-element group 192: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_352_Update/word_access_complete/word_0/ca
      -- 
    ca_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_352_store_0_ack_1, ack => initInputs_CP_117_elements(192)); -- 
    -- CP-element group 193:  transition  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	186 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	190 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_43/assign_stmt_344_to_assign_stmt_354/ptr_deref_343_ptr_deref_352_delay
      -- 
    -- Element group initInputs_CP_117_elements(193) is a control-delay.
    cp_element_193_delay: control_delay_element  generic map(name => " 193_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(186), ack => initInputs_CP_117_elements(193), clk => clk, reset =>reset);
    -- CP-element group 194:  transition  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	23 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (4) 
      -- CP-element group 194: 	 branch_block_stmt_43/assign_stmt_359/$entry
      -- CP-element group 194: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Sample/rr
      -- 
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(194), ack => RPIPE_rate_in_358_inst_req_0); -- 
    initInputs_CP_117_elements(194) <= initInputs_CP_117_elements(23);
    -- CP-element group 195:  transition  input  output  no-bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_update_start_
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Update/cr
      -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rate_in_358_inst_ack_0, ack => initInputs_CP_117_elements(195)); -- 
    cr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(195), ack => RPIPE_rate_in_358_inst_req_1); -- 
    -- CP-element group 196:  transition  input  no-bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	24 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_43/assign_stmt_359/$exit
      -- CP-element group 196: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_43/assign_stmt_359/RPIPE_rate_in_358_Update/ca
      -- 
    ca_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rate_in_358_inst_ack_1, ack => initInputs_CP_117_elements(196)); -- 
    -- CP-element group 197:  join  fork  transition  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	24 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	200 
    -- CP-element group 197: 	202 
    -- CP-element group 197: 	203 
    -- CP-element group 197: 	205 
    -- CP-element group 197:  members (59) 
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_update_start_
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_word_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_root_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_address_resized
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_addr_resize/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_addr_resize/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_addr_resize/base_resize_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_addr_resize/base_resize_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_plus_offset/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_plus_offset/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_plus_offset/sum_rename_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_base_plus_offset/sum_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_word_addrgen/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_word_addrgen/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_word_addrgen/root_register_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_word_addrgen/root_register_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/ptr_deref_361_Split/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/ptr_deref_361_Split/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/ptr_deref_361_Split/split_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/ptr_deref_361_Split/split_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/word_0/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/word_0/rr
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/word_0/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/word_0/cr
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_update_start_
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_word_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_root_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_address_resized
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_addr_resize/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_addr_resize/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_addr_resize/base_resize_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_addr_resize/base_resize_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_plus_offset/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_plus_offset/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_plus_offset/sum_rename_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_base_plus_offset/sum_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_word_addrgen/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_word_addrgen/$exit
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_word_addrgen/root_register_req
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_word_addrgen/root_register_ack
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/word_0/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/word_0/cr
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_update_start_
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_word_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_root_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/word_0/$entry
      -- CP-element group 197: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/word_0/cr
      -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(197), ack => ptr_deref_361_store_0_req_1); -- 
    rr_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(197), ack => ptr_deref_361_store_0_req_0); -- 
    cr_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(197), ack => ptr_deref_366_load_0_req_1); -- 
    cr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(197), ack => STORE_rate_368_store_0_req_1); -- 
    initInputs_CP_117_elements(197) <= initInputs_CP_117_elements(24);
    -- CP-element group 198:  transition  input  no-bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	206 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/$exit
      -- CP-element group 198: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/word_0/$exit
      -- CP-element group 198: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Sample/word_access_start/word_0/ra
      -- 
    ra_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_361_store_0_ack_0, ack => initInputs_CP_117_elements(198)); -- 
    -- CP-element group 199:  transition  input  no-bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	207 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/$exit
      -- CP-element group 199: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/word_0/$exit
      -- CP-element group 199: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_Update/word_access_complete/word_0/ca
      -- 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_361_store_0_ack_1, ack => initInputs_CP_117_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	197 
    -- CP-element group 200: 	206 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (5) 
      -- CP-element group 200: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/$entry
      -- CP-element group 200: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/word_0/$entry
      -- CP-element group 200: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/word_0/rr
      -- 
    rr_2240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(200), ack => ptr_deref_366_load_0_req_0); -- 
    initInputs_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(197) & initInputs_CP_117_elements(206);
      gj_initInputs_cp_element_group_200 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  no-bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (5) 
      -- CP-element group 201: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/$exit
      -- CP-element group 201: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/word_0/$exit
      -- CP-element group 201: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Sample/word_access_start/word_0/ra
      -- 
    ra_2241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_366_load_0_ack_0, ack => initInputs_CP_117_elements(201)); -- 
    -- CP-element group 202:  transition  input  no-bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (9) 
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/$exit
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/word_0/$exit
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/word_access_complete/word_0/ca
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/ptr_deref_366_Merge/$entry
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/ptr_deref_366_Merge/$exit
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/ptr_deref_366_Merge/merge_req
      -- CP-element group 202: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_366_Update/ptr_deref_366_Merge/merge_ack
      -- 
    ca_2252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_366_load_0_ack_1, ack => initInputs_CP_117_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	197 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/STORE_rate_368_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/STORE_rate_368_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/STORE_rate_368_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/STORE_rate_368_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/word_0/rr
      -- 
    rr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_117_elements(203), ack => STORE_rate_368_store_0_req_0); -- 
    initInputs_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(197) & initInputs_CP_117_elements(202);
      gj_initInputs_cp_element_group_203 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  no-bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Sample/word_access_start/word_0/ra
      -- 
    ra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_rate_368_store_0_ack_0, ack => initInputs_CP_117_elements(204)); -- 
    -- CP-element group 205:  transition  input  no-bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	197 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/STORE_rate_368_Update/word_access_complete/word_0/ca
      -- 
    ca_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_rate_368_store_0_ack_1, ack => initInputs_CP_117_elements(205)); -- 
    -- CP-element group 206:  transition  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	198 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	200 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/ptr_deref_361_ptr_deref_366_delay
      -- 
    -- Element group initInputs_CP_117_elements(206) is a control-delay.
    cp_element_206_delay: control_delay_element  generic map(name => " 206_delay", delay_value => 1)  port map(req => initInputs_CP_117_elements(198), ack => initInputs_CP_117_elements(206), clk => clk, reset =>reset);
    -- CP-element group 207:  join  transition  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	199 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	25 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_43/assign_stmt_363_to_assign_stmt_370/$exit
      -- 
    initInputs_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_117_elements(199) & initInputs_CP_117_elements(205);
      gj_initInputs_cp_element_group_207 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_117_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	6 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_43/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_43/bb_0_bb_1_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(208) <= initInputs_CP_117_elements(6);
    -- CP-element group 209:  transition  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	13 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_43/bb_3_bb_1_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_43/bb_3_bb_1_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(209) <= initInputs_CP_117_elements(13);
    -- CP-element group 210:  merge  place  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_43/merge_stmt_108_PhiReqMerge
      -- 
    initInputs_CP_117_elements(210) <= OrReduce(initInputs_CP_117_elements(208) & initInputs_CP_117_elements(209));
    -- CP-element group 211:  transition  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	7 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_43/merge_stmt_108_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_43/merge_stmt_108_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_43/merge_stmt_108_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(211) <= initInputs_CP_117_elements(210);
    -- CP-element group 212:  transition  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	72 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_43/bb_1_bb_2_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_43/bb_1_bb_2_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(212) <= initInputs_CP_117_elements(72);
    -- CP-element group 213:  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_43/merge_stmt_134_PhiReqMerge
      -- 
    initInputs_CP_117_elements(213) <= initInputs_CP_117_elements(212);
    -- CP-element group 214:  transition  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	9 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_43/merge_stmt_134_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_43/merge_stmt_134_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_43/merge_stmt_134_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(214) <= initInputs_CP_117_elements(213);
    -- CP-element group 215:  transition  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	11 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_43/bb_2_bb_3_PhiReq/$entry
      -- CP-element group 215: 	 branch_block_stmt_43/bb_2_bb_3_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(215) <= initInputs_CP_117_elements(11);
    -- CP-element group 216:  place  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 branch_block_stmt_43/merge_stmt_165_PhiReqMerge
      -- 
    initInputs_CP_117_elements(216) <= initInputs_CP_117_elements(215);
    -- CP-element group 217:  transition  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	12 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_43/merge_stmt_165_PhiAck/$entry
      -- CP-element group 217: 	 branch_block_stmt_43/merge_stmt_165_PhiAck/$exit
      -- CP-element group 217: 	 branch_block_stmt_43/merge_stmt_165_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(217) <= initInputs_CP_117_elements(216);
    -- CP-element group 218:  transition  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	73 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_43/bb_1_bb_4_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_43/bb_1_bb_4_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(218) <= initInputs_CP_117_elements(73);
    -- CP-element group 219:  place  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_43/merge_stmt_181_PhiReqMerge
      -- 
    initInputs_CP_117_elements(219) <= initInputs_CP_117_elements(218);
    -- CP-element group 220:  transition  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	14 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_43/merge_stmt_181_PhiAck/$entry
      -- CP-element group 220: 	 branch_block_stmt_43/merge_stmt_181_PhiAck/$exit
      -- CP-element group 220: 	 branch_block_stmt_43/merge_stmt_181_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(220) <= initInputs_CP_117_elements(219);
    -- CP-element group 221:  transition  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	15 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_43/bb_4_bb_5_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_43/bb_4_bb_5_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(221) <= initInputs_CP_117_elements(15);
    -- CP-element group 222:  transition  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	22 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_43/bb_7_bb_5_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_43/bb_7_bb_5_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(222) <= initInputs_CP_117_elements(22);
    -- CP-element group 223:  merge  place  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_43/merge_stmt_268_PhiReqMerge
      -- 
    initInputs_CP_117_elements(223) <= OrReduce(initInputs_CP_117_elements(221) & initInputs_CP_117_elements(222));
    -- CP-element group 224:  transition  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	16 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/$entry
      -- CP-element group 224: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/$exit
      -- CP-element group 224: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(224) <= initInputs_CP_117_elements(223);
    -- CP-element group 225:  transition  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	157 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_43/bb_5_bb_6_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_43/bb_5_bb_6_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(225) <= initInputs_CP_117_elements(157);
    -- CP-element group 226:  place  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_43/merge_stmt_298_PhiReqMerge
      -- 
    initInputs_CP_117_elements(226) <= initInputs_CP_117_elements(225);
    -- CP-element group 227:  transition  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	18 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_43/merge_stmt_298_PhiAck/$entry
      -- CP-element group 227: 	 branch_block_stmt_43/merge_stmt_298_PhiAck/$exit
      -- CP-element group 227: 	 branch_block_stmt_43/merge_stmt_298_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(227) <= initInputs_CP_117_elements(226);
    -- CP-element group 228:  transition  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	20 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_43/bb_6_bb_7_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_43/bb_6_bb_7_PhiReq/$exit
      -- 
    initInputs_CP_117_elements(228) <= initInputs_CP_117_elements(20);
    -- CP-element group 229:  place  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (1) 
      -- CP-element group 229: 	 branch_block_stmt_43/merge_stmt_340_PhiReqMerge
      -- 
    initInputs_CP_117_elements(229) <= initInputs_CP_117_elements(228);
    -- CP-element group 230:  transition  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	21 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_43/merge_stmt_340_PhiAck/dummy
      -- CP-element group 230: 	 branch_block_stmt_43/merge_stmt_340_PhiAck/$exit
      -- CP-element group 230: 	 branch_block_stmt_43/merge_stmt_340_PhiAck/$entry
      -- 
    initInputs_CP_117_elements(230) <= initInputs_CP_117_elements(229);
    -- CP-element group 231:  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	158 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_43/bb_5_bb_8_PhiReq/$exit
      -- CP-element group 231: 	 branch_block_stmt_43/bb_5_bb_8_PhiReq/$entry
      -- 
    initInputs_CP_117_elements(231) <= initInputs_CP_117_elements(158);
    -- CP-element group 232:  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_43/merge_stmt_356_PhiReqMerge
      -- 
    initInputs_CP_117_elements(232) <= initInputs_CP_117_elements(231);
    -- CP-element group 233:  transition  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	23 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_43/merge_stmt_356_PhiAck/dummy
      -- CP-element group 233: 	 branch_block_stmt_43/merge_stmt_356_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_43/merge_stmt_356_PhiAck/$entry
      -- 
    initInputs_CP_117_elements(233) <= initInputs_CP_117_elements(232);
    -- CP-element group 234:  transition  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	25 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_43/return___PhiReq/$entry
      -- CP-element group 234: 	 branch_block_stmt_43/return___PhiReq/$exit
      -- 
    initInputs_CP_117_elements(234) <= initInputs_CP_117_elements(25);
    -- CP-element group 235:  place  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (1) 
      -- CP-element group 235: 	 branch_block_stmt_43/merge_stmt_372_PhiReqMerge
      -- 
    initInputs_CP_117_elements(235) <= initInputs_CP_117_elements(234);
    -- CP-element group 236:  transition  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	26 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_43/merge_stmt_372_PhiAck/$entry
      -- CP-element group 236: 	 branch_block_stmt_43/merge_stmt_372_PhiAck/$exit
      -- CP-element group 236: 	 branch_block_stmt_43/merge_stmt_372_PhiAck/dummy
      -- 
    initInputs_CP_117_elements(236) <= initInputs_CP_117_elements(235);
    -- CP-element group 237:  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	26 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 $exit
      -- CP-element group 237: 	 branch_block_stmt_43/$exit
      -- 
    initInputs_CP_117_elements(237) <= initInputs_CP_117_elements(26);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_61 : std_logic_vector(31 downto 0);
    signal R_iNsTr_21_156_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_21_156_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_63_331_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_63_331_scaled : std_logic_vector(9 downto 0);
    signal Rate_73 : std_logic_vector(31 downto 0);
    signal SNR_57 : std_logic_vector(31 downto 0);
    signal STORE_ebbyNo_99_data_0 : std_logic_vector(31 downto 0);
    signal STORE_ebbyNo_99_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_maxNitr_85_data_0 : std_logic_vector(15 downto 0);
    signal STORE_maxNitr_85_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ncol_ind_218_data_0 : std_logic_vector(15 downto 0);
    signal STORE_ncol_ind_218_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ncols_205_data_0 : std_logic_vector(15 downto 0);
    signal STORE_ncols_205_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_nrows_192_data_0 : std_logic_vector(15 downto 0);
    signal STORE_nrows_192_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_rate_368_data_0 : std_logic_vector(31 downto 0);
    signal STORE_rate_368_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_157_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_157_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_157_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_157_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_332_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_332_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_332_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_332_root_address : std_logic_vector(9 downto 0);
    signal iNsTr_12_112 : std_logic_vector(15 downto 0);
    signal iNsTr_13_117 : std_logic_vector(31 downto 0);
    signal iNsTr_14_127 : std_logic_vector(0 downto 0);
    signal iNsTr_17_137 : std_logic_vector(15 downto 0);
    signal iNsTr_19_145 : std_logic_vector(15 downto 0);
    signal iNsTr_1_76 : std_logic_vector(15 downto 0);
    signal iNsTr_20_149 : std_logic_vector(15 downto 0);
    signal iNsTr_21_154 : std_logic_vector(63 downto 0);
    signal iNsTr_22_159 : std_logic_vector(31 downto 0);
    signal iNsTr_25_187 : std_logic_vector(31 downto 0);
    signal iNsTr_26_191 : std_logic_vector(15 downto 0);
    signal iNsTr_28_200 : std_logic_vector(31 downto 0);
    signal iNsTr_29_204 : std_logic_vector(15 downto 0);
    signal iNsTr_31_213 : std_logic_vector(31 downto 0);
    signal iNsTr_32_217 : std_logic_vector(15 downto 0);
    signal iNsTr_34_226 : std_logic_vector(31 downto 0);
    signal iNsTr_35_230 : std_logic_vector(15 downto 0);
    signal iNsTr_36_234 : std_logic_vector(31 downto 0);
    signal iNsTr_37_240 : std_logic_vector(31 downto 0);
    signal iNsTr_38_244 : std_logic_vector(15 downto 0);
    signal iNsTr_39_248 : std_logic_vector(31 downto 0);
    signal iNsTr_3_84 : std_logic_vector(15 downto 0);
    signal iNsTr_40_253 : std_logic_vector(31 downto 0);
    signal iNsTr_41_257 : std_logic_vector(15 downto 0);
    signal iNsTr_45_169 : std_logic_vector(15 downto 0);
    signal iNsTr_46_175 : std_logic_vector(15 downto 0);
    signal iNsTr_49_272 : std_logic_vector(15 downto 0);
    signal iNsTr_50_276 : std_logic_vector(31 downto 0);
    signal iNsTr_51_280 : std_logic_vector(15 downto 0);
    signal iNsTr_52_284 : std_logic_vector(31 downto 0);
    signal iNsTr_53_291 : std_logic_vector(0 downto 0);
    signal iNsTr_57_301 : std_logic_vector(15 downto 0);
    signal iNsTr_59_309 : std_logic_vector(15 downto 0);
    signal iNsTr_60_313 : std_logic_vector(15 downto 0);
    signal iNsTr_61_317 : std_logic_vector(31 downto 0);
    signal iNsTr_62_323 : std_logic_vector(31 downto 0);
    signal iNsTr_63_329 : std_logic_vector(63 downto 0);
    signal iNsTr_64_334 : std_logic_vector(31 downto 0);
    signal iNsTr_68_359 : std_logic_vector(31 downto 0);
    signal iNsTr_6_90 : std_logic_vector(31 downto 0);
    signal iNsTr_70_367 : std_logic_vector(31 downto 0);
    signal iNsTr_73_344 : std_logic_vector(15 downto 0);
    signal iNsTr_74_350 : std_logic_vector(15 downto 0);
    signal iNsTr_8_98 : std_logic_vector(31 downto 0);
    signal nitr_53 : std_logic_vector(31 downto 0);
    signal ptr_deref_103_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_103_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_103_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_103_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_103_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_103_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_111_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_111_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_111_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_111_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_111_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_139_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_139_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_139_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_139_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_139_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_139_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_144_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_144_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_144_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_144_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_144_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_148_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_148_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_148_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_148_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_148_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_161_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_161_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_161_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_161_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_161_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_161_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_168_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_168_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_168_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_168_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_168_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_177_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_177_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_177_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_177_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_177_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_177_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_190_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_190_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_190_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_190_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_190_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_203_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_203_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_203_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_203_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_203_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_216_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_216_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_216_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_216_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_216_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_229_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_229_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_229_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_229_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_229_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_243_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_243_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_243_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_243_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_243_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_259_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_259_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_259_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_259_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_259_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_259_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_263_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_263_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_263_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_271_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_271_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_271_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_271_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_271_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_279_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_279_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_279_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_279_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_279_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_303_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_303_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_303_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_303_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_303_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_303_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_308_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_308_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_308_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_308_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_308_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_312_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_312_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_312_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_312_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_312_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_336_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_336_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_336_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_336_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_336_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_336_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_343_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_343_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_343_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_352_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_352_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_352_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_352_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_352_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_352_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_361_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_361_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_361_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_361_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_361_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_361_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_366_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_366_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_366_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_366_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_366_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_78_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_78_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_78_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_78_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_78_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_78_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_83_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_83_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_83_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_83_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_83_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_92_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_92_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_92_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_92_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_92_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_92_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_97_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_97_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_97_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_97_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_97_word_offset_0 : std_logic_vector(0 downto 0);
    signal range_69 : std_logic_vector(31 downto 0);
    signal type_cast_105_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_121_wire : std_logic_vector(31 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_173_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_265_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_287_wire : std_logic_vector(31 downto 0);
    signal type_cast_289_wire : std_logic_vector(31 downto 0);
    signal type_cast_321_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_327_wire : std_logic_vector(63 downto 0);
    signal type_cast_348_wire_constant : std_logic_vector(15 downto 0);
    signal val_65 : std_logic_vector(31 downto 0);
    signal xxinitInputsxxbodyxxI_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinitInputsxxbodyxxRate_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinitInputsxxbodyxxSNR_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinitInputsxxbodyxxnitr_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinitInputsxxbodyxxrange_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinitInputsxxbodyxxval_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    I_61 <= "00000000000000000000000000000000";
    Rate_73 <= "00000000000000000000000000000000";
    SNR_57 <= "00000000000000000000000000000000";
    STORE_ebbyNo_99_word_address_0 <= "0";
    STORE_maxNitr_85_word_address_0 <= "0";
    STORE_ncol_ind_218_word_address_0 <= "0";
    STORE_ncols_205_word_address_0 <= "0";
    STORE_nrows_192_word_address_0 <= "0";
    STORE_rate_368_word_address_0 <= "0";
    array_obj_ref_157_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_157_resized_base_address <= "0000000000";
    array_obj_ref_332_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_332_resized_base_address <= "0000000000";
    iNsTr_25_187 <= "00000000000000000000000000000000";
    iNsTr_28_200 <= "00000000000000000000000000000001";
    iNsTr_31_213 <= "00000000000000000000000000000010";
    iNsTr_34_226 <= "00000000000000000000000000000010";
    iNsTr_37_240 <= "00000000000000000000000000000000";
    nitr_53 <= "00000000000000000000000000000000";
    ptr_deref_103_word_offset_0 <= "0";
    ptr_deref_111_word_offset_0 <= "0";
    ptr_deref_139_word_offset_0 <= "0";
    ptr_deref_144_word_offset_0 <= "0";
    ptr_deref_148_word_offset_0 <= "0";
    ptr_deref_161_word_offset_0 <= "0000000000";
    ptr_deref_168_word_offset_0 <= "0";
    ptr_deref_177_word_offset_0 <= "0";
    ptr_deref_190_word_offset_0 <= "0000000000";
    ptr_deref_203_word_offset_0 <= "0000000000";
    ptr_deref_216_word_offset_0 <= "0000000000";
    ptr_deref_229_word_offset_0 <= "0000000000";
    ptr_deref_243_word_offset_0 <= "0000000000";
    ptr_deref_259_word_offset_0 <= "0";
    ptr_deref_263_word_offset_0 <= "0";
    ptr_deref_271_word_offset_0 <= "0";
    ptr_deref_279_word_offset_0 <= "0";
    ptr_deref_303_word_offset_0 <= "0";
    ptr_deref_308_word_offset_0 <= "0";
    ptr_deref_312_word_offset_0 <= "0";
    ptr_deref_336_word_offset_0 <= "0000000000";
    ptr_deref_343_word_offset_0 <= "0";
    ptr_deref_352_word_offset_0 <= "0";
    ptr_deref_361_word_offset_0 <= "0";
    ptr_deref_366_word_offset_0 <= "0";
    ptr_deref_78_word_offset_0 <= "0";
    ptr_deref_83_word_offset_0 <= "0";
    ptr_deref_92_word_offset_0 <= "0";
    ptr_deref_97_word_offset_0 <= "0";
    range_69 <= "00000000000000000000000000000000";
    type_cast_105_wire_constant <= "0000000000000000";
    type_cast_124_wire_constant <= "00000000000000000000000000000011";
    type_cast_173_wire_constant <= "0000000000000001";
    type_cast_265_wire_constant <= "0000000000000000";
    type_cast_321_wire_constant <= "00000000000000000000000000000011";
    type_cast_348_wire_constant <= "0000000000000001";
    val_65 <= "00000000000000000000000000000000";
    xxinitInputsxxbodyxxI_alloc_base_address <= "0";
    xxinitInputsxxbodyxxRate_alloc_base_address <= "0";
    xxinitInputsxxbodyxxSNR_alloc_base_address <= "0";
    xxinitInputsxxbodyxxnitr_alloc_base_address <= "0";
    xxinitInputsxxbodyxxrange_alloc_base_address <= "0";
    xxinitInputsxxbodyxxval_alloc_base_address <= "0";
    addr_of_158_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_158_final_reg_req_0;
      addr_of_158_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_158_final_reg_req_1;
      addr_of_158_final_reg_ack_1<= rack(0);
      addr_of_158_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_158_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_157_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_22_159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_333_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_333_final_reg_req_0;
      addr_of_333_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_333_final_reg_req_1;
      addr_of_333_final_reg_ack_1<= rack(0);
      addr_of_333_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_333_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_332_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_64_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_116_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_116_inst_req_0;
      type_cast_116_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_116_inst_req_1;
      type_cast_116_inst_ack_1<= rack(0);
      type_cast_116_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_116_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_12_112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_13_117,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_121_inst
    process(iNsTr_13_117) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_13_117(31 downto 0);
      type_cast_121_wire <= tmp_var; -- 
    end process;
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_20_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_21_154,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_233_inst_req_0;
      type_cast_233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_233_inst_req_1;
      type_cast_233_inst_ack_1<= rack(0);
      type_cast_233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_36_234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_247_inst_req_0;
      type_cast_247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_247_inst_req_1;
      type_cast_247_inst_ack_1<= rack(0);
      type_cast_247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_38_244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_256_inst_req_0;
      type_cast_256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_256_inst_req_1;
      type_cast_256_inst_ack_1<= rack(0);
      type_cast_256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_40_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_41_257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_275_inst_req_0;
      type_cast_275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_275_inst_req_1;
      type_cast_275_inst_ack_1<= rack(0);
      type_cast_275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_49_272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_50_276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_283_inst_req_0;
      type_cast_283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_283_inst_req_1;
      type_cast_283_inst_ack_1<= rack(0);
      type_cast_283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_51_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_287_inst
    process(iNsTr_50_276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_50_276(31 downto 0);
      type_cast_287_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_289_inst
    process(iNsTr_52_284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_52_284(31 downto 0);
      type_cast_289_wire <= tmp_var; -- 
    end process;
    type_cast_316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_316_inst_req_0;
      type_cast_316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_316_inst_req_1;
      type_cast_316_inst_ack_1<= rack(0);
      type_cast_316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_60_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_61_317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_328_inst_req_0;
      type_cast_328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_328_inst_req_1;
      type_cast_328_inst_ack_1<= rack(0);
      type_cast_328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_327_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_63_329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_ebbyNo_99_gather_scatter
    process(iNsTr_8_98) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_98;
      ov(31 downto 0) := iv;
      STORE_ebbyNo_99_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_maxNitr_85_gather_scatter
    process(iNsTr_3_84) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_84;
      ov(15 downto 0) := iv;
      STORE_maxNitr_85_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_ncol_ind_218_gather_scatter
    process(iNsTr_32_217) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_217;
      ov(15 downto 0) := iv;
      STORE_ncol_ind_218_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_ncols_205_gather_scatter
    process(iNsTr_29_204) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_204;
      ov(15 downto 0) := iv;
      STORE_ncols_205_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_nrows_192_gather_scatter
    process(iNsTr_26_191) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_191;
      ov(15 downto 0) := iv;
      STORE_nrows_192_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_rate_368_gather_scatter
    process(iNsTr_70_367) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_70_367;
      ov(31 downto 0) := iv;
      STORE_rate_368_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_157_index_0_rename
    process(R_iNsTr_21_156_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_21_156_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_21_156_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_157_index_0_resize
    process(iNsTr_21_154) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_154;
      ov := iv(9 downto 0);
      R_iNsTr_21_156_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_157_index_offset
    process(R_iNsTr_21_156_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_21_156_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_157_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_157_root_address_inst
    process(array_obj_ref_157_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_157_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_157_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_332_index_0_rename
    process(R_iNsTr_63_331_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_63_331_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_63_331_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_332_index_0_resize
    process(iNsTr_63_329) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_63_329;
      ov := iv(9 downto 0);
      R_iNsTr_63_331_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_332_index_offset
    process(R_iNsTr_63_331_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_63_331_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_332_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_332_root_address_inst
    process(array_obj_ref_332_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_332_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_332_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_103_addr_0
    process(ptr_deref_103_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_103_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_103_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_103_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_103_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_103_gather_scatter
    process(type_cast_105_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_105_wire_constant;
      ov(15 downto 0) := iv;
      ptr_deref_103_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_103_root_address_inst
    process(ptr_deref_103_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_103_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_103_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_111_addr_0
    process(ptr_deref_111_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_111_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_111_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_111_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_111_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_111_gather_scatter
    process(ptr_deref_111_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_111_data_0;
      ov(15 downto 0) := iv;
      iNsTr_12_112 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_111_root_address_inst
    process(ptr_deref_111_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_111_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_111_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_addr_0
    process(ptr_deref_139_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_139_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_base_resize
    process(val_65) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_65;
      ov := iv(0 downto 0);
      ptr_deref_139_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_gather_scatter
    process(iNsTr_17_137) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_137;
      ov(15 downto 0) := iv;
      ptr_deref_139_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_root_address_inst
    process(ptr_deref_139_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_139_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_144_addr_0
    process(ptr_deref_144_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_144_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_144_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_144_base_resize
    process(val_65) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_65;
      ov := iv(0 downto 0);
      ptr_deref_144_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_144_gather_scatter
    process(ptr_deref_144_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_144_data_0;
      ov(15 downto 0) := iv;
      iNsTr_19_145 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_144_root_address_inst
    process(ptr_deref_144_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_144_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_144_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_addr_0
    process(ptr_deref_148_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_148_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_148_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_gather_scatter
    process(ptr_deref_148_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_data_0;
      ov(15 downto 0) := iv;
      iNsTr_20_149 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_root_address_inst
    process(ptr_deref_148_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_148_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_161_addr_0
    process(ptr_deref_161_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_161_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_161_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_161_base_resize
    process(iNsTr_22_159) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_159;
      ov := iv(9 downto 0);
      ptr_deref_161_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_161_gather_scatter
    process(iNsTr_19_145) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_145;
      ov(15 downto 0) := iv;
      ptr_deref_161_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_161_root_address_inst
    process(ptr_deref_161_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_161_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_161_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_168_addr_0
    process(ptr_deref_168_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_168_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_168_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_168_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_168_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_168_gather_scatter
    process(ptr_deref_168_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_168_data_0;
      ov(15 downto 0) := iv;
      iNsTr_45_169 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_168_root_address_inst
    process(ptr_deref_168_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_168_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_168_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_177_addr_0
    process(ptr_deref_177_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_177_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_177_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_177_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_177_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_177_gather_scatter
    process(iNsTr_46_175) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_175;
      ov(15 downto 0) := iv;
      ptr_deref_177_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_177_root_address_inst
    process(ptr_deref_177_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_177_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_177_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_190_addr_0
    process(ptr_deref_190_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_190_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_190_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_190_base_resize
    process(iNsTr_25_187) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_187;
      ov := iv(9 downto 0);
      ptr_deref_190_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_190_gather_scatter
    process(ptr_deref_190_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_190_data_0;
      ov(15 downto 0) := iv;
      iNsTr_26_191 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_190_root_address_inst
    process(ptr_deref_190_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_190_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_190_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_203_addr_0
    process(ptr_deref_203_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_203_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_203_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_203_base_resize
    process(iNsTr_28_200) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_28_200;
      ov := iv(9 downto 0);
      ptr_deref_203_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_203_gather_scatter
    process(ptr_deref_203_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_203_data_0;
      ov(15 downto 0) := iv;
      iNsTr_29_204 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_203_root_address_inst
    process(ptr_deref_203_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_203_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_203_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_addr_0
    process(ptr_deref_216_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_216_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_216_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_base_resize
    process(iNsTr_31_213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_31_213;
      ov := iv(9 downto 0);
      ptr_deref_216_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_gather_scatter
    process(ptr_deref_216_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_216_data_0;
      ov(15 downto 0) := iv;
      iNsTr_32_217 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_root_address_inst
    process(ptr_deref_216_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_216_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_216_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_229_addr_0
    process(ptr_deref_229_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_229_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_229_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_229_base_resize
    process(iNsTr_34_226) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_226;
      ov := iv(9 downto 0);
      ptr_deref_229_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_229_gather_scatter
    process(ptr_deref_229_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_229_data_0;
      ov(15 downto 0) := iv;
      iNsTr_35_230 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_229_root_address_inst
    process(ptr_deref_229_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_229_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_229_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_243_addr_0
    process(ptr_deref_243_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_243_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_243_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_243_base_resize
    process(iNsTr_37_240) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_240;
      ov := iv(9 downto 0);
      ptr_deref_243_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_243_gather_scatter
    process(ptr_deref_243_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_243_data_0;
      ov(15 downto 0) := iv;
      iNsTr_38_244 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_243_root_address_inst
    process(ptr_deref_243_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_243_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_243_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_259_addr_0
    process(ptr_deref_259_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_259_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_259_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_259_base_resize
    process(range_69) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := range_69;
      ov := iv(0 downto 0);
      ptr_deref_259_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_259_gather_scatter
    process(iNsTr_41_257) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_41_257;
      ov(15 downto 0) := iv;
      ptr_deref_259_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_259_root_address_inst
    process(ptr_deref_259_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_259_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_259_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_addr_0
    process(ptr_deref_263_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_263_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_263_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_gather_scatter
    process(type_cast_265_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_265_wire_constant;
      ov(15 downto 0) := iv;
      ptr_deref_263_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_root_address_inst
    process(ptr_deref_263_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_263_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_271_addr_0
    process(ptr_deref_271_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_271_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_271_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_271_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_271_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_271_gather_scatter
    process(ptr_deref_271_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_271_data_0;
      ov(15 downto 0) := iv;
      iNsTr_49_272 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_271_root_address_inst
    process(ptr_deref_271_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_271_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_271_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_addr_0
    process(ptr_deref_279_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_279_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_279_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_base_resize
    process(range_69) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := range_69;
      ov := iv(0 downto 0);
      ptr_deref_279_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_gather_scatter
    process(ptr_deref_279_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_279_data_0;
      ov(15 downto 0) := iv;
      iNsTr_51_280 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_279_root_address_inst
    process(ptr_deref_279_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_279_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_279_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_addr_0
    process(ptr_deref_303_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_303_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_base_resize
    process(val_65) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_65;
      ov := iv(0 downto 0);
      ptr_deref_303_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_gather_scatter
    process(iNsTr_57_301) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_57_301;
      ov(15 downto 0) := iv;
      ptr_deref_303_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_root_address_inst
    process(ptr_deref_303_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_303_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_308_addr_0
    process(ptr_deref_308_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_308_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_308_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_308_base_resize
    process(val_65) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_65;
      ov := iv(0 downto 0);
      ptr_deref_308_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_308_gather_scatter
    process(ptr_deref_308_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_308_data_0;
      ov(15 downto 0) := iv;
      iNsTr_59_309 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_308_root_address_inst
    process(ptr_deref_308_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_308_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_308_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_312_addr_0
    process(ptr_deref_312_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_312_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_312_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_312_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_312_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_312_gather_scatter
    process(ptr_deref_312_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_312_data_0;
      ov(15 downto 0) := iv;
      iNsTr_60_313 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_312_root_address_inst
    process(ptr_deref_312_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_312_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_312_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_336_addr_0
    process(ptr_deref_336_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_336_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_336_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_336_base_resize
    process(iNsTr_64_334) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_64_334;
      ov := iv(9 downto 0);
      ptr_deref_336_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_336_gather_scatter
    process(iNsTr_59_309) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_59_309;
      ov(15 downto 0) := iv;
      ptr_deref_336_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_336_root_address_inst
    process(ptr_deref_336_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_336_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_336_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_addr_0
    process(ptr_deref_343_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_343_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_343_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_gather_scatter
    process(ptr_deref_343_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_data_0;
      ov(15 downto 0) := iv;
      iNsTr_73_344 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_root_address_inst
    process(ptr_deref_343_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_343_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_352_addr_0
    process(ptr_deref_352_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_352_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_352_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_352_base_resize
    process(I_61) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_61;
      ov := iv(0 downto 0);
      ptr_deref_352_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_352_gather_scatter
    process(iNsTr_74_350) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_74_350;
      ov(15 downto 0) := iv;
      ptr_deref_352_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_352_root_address_inst
    process(ptr_deref_352_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_352_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_352_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_361_addr_0
    process(ptr_deref_361_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_361_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_361_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_361_base_resize
    process(Rate_73) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Rate_73;
      ov := iv(0 downto 0);
      ptr_deref_361_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_361_gather_scatter
    process(iNsTr_68_359) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_68_359;
      ov(31 downto 0) := iv;
      ptr_deref_361_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_361_root_address_inst
    process(ptr_deref_361_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_361_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_361_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_366_addr_0
    process(ptr_deref_366_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_366_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_366_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_366_base_resize
    process(Rate_73) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Rate_73;
      ov := iv(0 downto 0);
      ptr_deref_366_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_366_gather_scatter
    process(ptr_deref_366_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_366_data_0;
      ov(31 downto 0) := iv;
      iNsTr_70_367 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_366_root_address_inst
    process(ptr_deref_366_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_366_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_366_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_78_addr_0
    process(ptr_deref_78_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_78_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_78_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_78_base_resize
    process(nitr_53) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := nitr_53;
      ov := iv(0 downto 0);
      ptr_deref_78_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_78_gather_scatter
    process(iNsTr_1_76) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_76;
      ov(15 downto 0) := iv;
      ptr_deref_78_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_78_root_address_inst
    process(ptr_deref_78_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_78_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_78_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_83_addr_0
    process(ptr_deref_83_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_83_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_83_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_83_base_resize
    process(nitr_53) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := nitr_53;
      ov := iv(0 downto 0);
      ptr_deref_83_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_83_gather_scatter
    process(ptr_deref_83_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_83_data_0;
      ov(15 downto 0) := iv;
      iNsTr_3_84 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_83_root_address_inst
    process(ptr_deref_83_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_83_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_83_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_92_addr_0
    process(ptr_deref_92_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_92_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_92_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_92_base_resize
    process(SNR_57) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := SNR_57;
      ov := iv(0 downto 0);
      ptr_deref_92_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_92_gather_scatter
    process(iNsTr_6_90) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_90;
      ov(31 downto 0) := iv;
      ptr_deref_92_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_92_root_address_inst
    process(ptr_deref_92_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_92_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_92_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_97_addr_0
    process(ptr_deref_97_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_97_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_97_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_97_base_resize
    process(SNR_57) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := SNR_57;
      ov := iv(0 downto 0);
      ptr_deref_97_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_97_gather_scatter
    process(ptr_deref_97_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_97_data_0;
      ov(31 downto 0) := iv;
      iNsTr_8_98 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_97_root_address_inst
    process(ptr_deref_97_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_97_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_97_root_address <= ov(0 downto 0);
      --
    end process;
    if_stmt_128_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_14_127;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_128_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_128_branch_req_0,
          ack0 => if_stmt_128_branch_ack_0,
          ack1 => if_stmt_128_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_292_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_53_291;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_292_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_292_branch_req_0,
          ack0 => if_stmt_292_branch_ack_0,
          ack1 => if_stmt_292_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u16_u16_174_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_45_169;
      iNsTr_46_175 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_174_inst_req_0;
      ADD_u16_u16_174_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_174_inst_req_1;
      ADD_u16_u16_174_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u16_u16_349_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_73_344;
      iNsTr_74_350 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_349_inst_req_0;
      ADD_u16_u16_349_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_349_inst_req_1;
      ADD_u16_u16_349_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u32_u32_252_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_36_234 & iNsTr_39_248;
      iNsTr_40_253 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_252_inst_req_0;
      ADD_u32_u32_252_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_252_inst_req_1;
      ADD_u32_u32_252_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u32_u32_322_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_61_317;
      iNsTr_62_323 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_322_inst_req_0;
      ADD_u32_u32_322_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_322_inst_req_1;
      ADD_u32_u32_322_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : SLT_i32_u1_125_inst 
    ApIntSlt_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_121_wire;
      iNsTr_14_127 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_125_inst_req_0;
      SLT_i32_u1_125_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_125_inst_req_1;
      SLT_i32_u1_125_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_4_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : SLT_i32_u1_290_inst 
    ApIntSlt_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_287_wire & type_cast_289_wire;
      iNsTr_53_291 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_290_inst_req_0;
      SLT_i32_u1_290_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_290_inst_req_1;
      SLT_i32_u1_290_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_5_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : type_cast_327_inst 
    ApIntToApIntSigned_group_6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_62_323;
      type_cast_327_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_327_inst_req_0;
      type_cast_327_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_327_inst_req_1;
      type_cast_327_inst_ack_1 <= ackR_unguarded(0);
      ApIntToApIntSigned_group_6_gI: SplitGuardInterface generic map(name => "ApIntToApIntSigned_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared load operator group (0) : ptr_deref_271_load_0 ptr_deref_343_load_0 ptr_deref_111_load_0 ptr_deref_148_load_0 ptr_deref_168_load_0 ptr_deref_312_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_271_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_343_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_111_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_148_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_168_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_312_load_0_req_0;
      ptr_deref_271_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_343_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_111_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_148_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_168_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_312_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_271_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_343_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_111_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_148_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_168_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_312_load_0_req_1;
      ptr_deref_271_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_343_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_111_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_148_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_168_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_312_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_271_word_address_0 & ptr_deref_343_word_address_0 & ptr_deref_111_word_address_0 & ptr_deref_148_word_address_0 & ptr_deref_168_word_address_0 & ptr_deref_312_word_address_0;
      ptr_deref_271_data_0 <= data_out(95 downto 80);
      ptr_deref_343_data_0 <= data_out(79 downto 64);
      ptr_deref_111_data_0 <= data_out(63 downto 48);
      ptr_deref_148_data_0 <= data_out(47 downto 32);
      ptr_deref_168_data_0 <= data_out(31 downto 16);
      ptr_deref_312_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(0),
          mack => memory_space_11_lr_ack(0),
          maddr => memory_space_11_lr_addr(0 downto 0),
          mtag => memory_space_11_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(0),
          mack => memory_space_11_lc_ack(0),
          mdata => memory_space_11_lc_data(15 downto 0),
          mtag => memory_space_11_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_308_load_0 ptr_deref_144_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_308_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_144_load_0_req_0;
      ptr_deref_308_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_144_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_308_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_144_load_0_req_1;
      ptr_deref_308_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_144_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_308_word_address_0 & ptr_deref_144_word_address_0;
      ptr_deref_308_data_0 <= data_out(31 downto 16);
      ptr_deref_144_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_12_lr_req(0),
          mack => memory_space_12_lr_ack(0),
          maddr => memory_space_12_lr_addr(0 downto 0),
          mtag => memory_space_12_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_12_lc_req(0),
          mack => memory_space_12_lc_ack(0),
          mdata => memory_space_12_lc_data(15 downto 0),
          mtag => memory_space_12_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_229_load_0 ptr_deref_243_load_0 ptr_deref_216_load_0 ptr_deref_203_load_0 ptr_deref_190_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(49 downto 0);
      signal data_out: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_229_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_243_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_216_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_203_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_190_load_0_req_0;
      ptr_deref_229_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_243_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_216_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_203_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_190_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_229_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_243_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_216_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_203_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_190_load_0_req_1;
      ptr_deref_229_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_243_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_216_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_203_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_190_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_229_word_address_0 & ptr_deref_243_word_address_0 & ptr_deref_216_word_address_0 & ptr_deref_203_word_address_0 & ptr_deref_190_word_address_0;
      ptr_deref_229_data_0 <= data_out(79 downto 64);
      ptr_deref_243_data_0 <= data_out(63 downto 48);
      ptr_deref_216_data_0 <= data_out(47 downto 32);
      ptr_deref_203_data_0 <= data_out(31 downto 16);
      ptr_deref_190_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 10,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(9 downto 0),
          mtag => memory_space_4_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(15 downto 0),
          mtag => memory_space_4_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_279_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_279_load_0_req_0;
      ptr_deref_279_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_279_load_0_req_1;
      ptr_deref_279_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_279_word_address_0;
      ptr_deref_279_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_13_lr_req(0),
          mack => memory_space_13_lr_ack(0),
          maddr => memory_space_13_lr_addr(0 downto 0),
          mtag => memory_space_13_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_13_lc_req(0),
          mack => memory_space_13_lc_ack(0),
          mdata => memory_space_13_lc_data(15 downto 0),
          mtag => memory_space_13_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_366_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_366_load_0_req_0;
      ptr_deref_366_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_366_load_0_req_1;
      ptr_deref_366_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_366_word_address_0;
      ptr_deref_366_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_14_lr_req(0),
          mack => memory_space_14_lr_ack(0),
          maddr => memory_space_14_lr_addr(0 downto 0),
          mtag => memory_space_14_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_14_lc_req(0),
          mack => memory_space_14_lc_ack(0),
          mdata => memory_space_14_lc_data(31 downto 0),
          mtag => memory_space_14_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_83_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_83_load_0_req_0;
      ptr_deref_83_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_83_load_0_req_1;
      ptr_deref_83_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_83_word_address_0;
      ptr_deref_83_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(0 downto 0),
          mtag => memory_space_9_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(15 downto 0),
          mtag => memory_space_9_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_97_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_97_load_0_req_0;
      ptr_deref_97_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_97_load_0_req_1;
      ptr_deref_97_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_97_word_address_0;
      ptr_deref_97_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(31 downto 0),
          mtag => memory_space_10_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared store operator group (0) : STORE_ebbyNo_99_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ebbyNo_99_store_0_req_0;
      STORE_ebbyNo_99_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ebbyNo_99_store_0_req_1;
      STORE_ebbyNo_99_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ebbyNo_99_word_address_0;
      data_in <= STORE_ebbyNo_99_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_maxNitr_85_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_maxNitr_85_store_0_req_0;
      STORE_maxNitr_85_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_maxNitr_85_store_0_req_1;
      STORE_maxNitr_85_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_maxNitr_85_word_address_0;
      data_in <= STORE_maxNitr_85_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(0 downto 0),
          mdata => memory_space_3_sr_data(15 downto 0),
          mtag => memory_space_3_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_ncol_ind_218_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ncol_ind_218_store_0_req_0;
      STORE_ncol_ind_218_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ncol_ind_218_store_0_req_1;
      STORE_ncol_ind_218_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ncol_ind_218_word_address_0;
      data_in <= STORE_ncol_ind_218_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(0 downto 0),
          mdata => memory_space_5_sr_data(15 downto 0),
          mtag => memory_space_5_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : STORE_ncols_205_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ncols_205_store_0_req_0;
      STORE_ncols_205_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ncols_205_store_0_req_1;
      STORE_ncols_205_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ncols_205_word_address_0;
      data_in <= STORE_ncols_205_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : STORE_nrows_192_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_nrows_192_store_0_req_0;
      STORE_nrows_192_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_nrows_192_store_0_req_1;
      STORE_nrows_192_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_nrows_192_word_address_0;
      data_in <= STORE_nrows_192_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : STORE_rate_368_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_rate_368_store_0_req_0;
      STORE_rate_368_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_rate_368_store_0_req_1;
      STORE_rate_368_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_rate_368_word_address_0;
      data_in <= STORE_rate_368_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(31 downto 0),
          mtag => memory_space_8_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_352_store_0 ptr_deref_263_store_0 ptr_deref_103_store_0 ptr_deref_177_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_352_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_263_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_103_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_177_store_0_req_0;
      ptr_deref_352_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_263_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_103_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_177_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_352_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_263_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_103_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_177_store_0_req_1;
      ptr_deref_352_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_263_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_103_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_177_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup6_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_352_word_address_0 & ptr_deref_263_word_address_0 & ptr_deref_103_word_address_0 & ptr_deref_177_word_address_0;
      data_in <= ptr_deref_352_data_0 & ptr_deref_263_data_0 & ptr_deref_103_data_0 & ptr_deref_177_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(0 downto 0),
          mdata => memory_space_11_sr_data(15 downto 0),
          mtag => memory_space_11_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_303_store_0 ptr_deref_139_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_303_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_139_store_0_req_0;
      ptr_deref_303_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_139_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_303_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_139_store_0_req_1;
      ptr_deref_303_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_139_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup7_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup7_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup7_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup7_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_303_word_address_0 & ptr_deref_139_word_address_0;
      data_in <= ptr_deref_303_data_0 & ptr_deref_139_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_12_sr_req(0),
          mack => memory_space_12_sr_ack(0),
          maddr => memory_space_12_sr_addr(0 downto 0),
          mdata => memory_space_12_sr_data(15 downto 0),
          mtag => memory_space_12_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_12_sc_req(0),
          mack => memory_space_12_sc_ack(0),
          mtag => memory_space_12_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : ptr_deref_336_store_0 ptr_deref_161_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(19 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_336_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_161_store_0_req_0;
      ptr_deref_336_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_161_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_336_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_161_store_0_req_1;
      ptr_deref_336_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_161_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup8_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup8_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup8_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup8_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup8_gI: SplitGuardInterface generic map(name => "StoreGroup8_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_336_word_address_0 & ptr_deref_161_word_address_0;
      data_in <= ptr_deref_336_data_0 & ptr_deref_161_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup8 Req ", addr_width => 10,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(9 downto 0),
          mdata => memory_space_4_sr_data(15 downto 0),
          mtag => memory_space_4_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup8 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared store operator group (9) : ptr_deref_259_store_0 
    StoreGroup9: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_259_store_0_req_0;
      ptr_deref_259_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_259_store_0_req_1;
      ptr_deref_259_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup9_gI: SplitGuardInterface generic map(name => "StoreGroup9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_259_word_address_0;
      data_in <= ptr_deref_259_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup9 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_13_sr_req(0),
          mack => memory_space_13_sr_ack(0),
          maddr => memory_space_13_sr_addr(0 downto 0),
          mdata => memory_space_13_sr_data(15 downto 0),
          mtag => memory_space_13_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup9 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_13_sc_req(0),
          mack => memory_space_13_sc_ack(0),
          mtag => memory_space_13_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 9
    -- shared store operator group (10) : ptr_deref_361_store_0 
    StoreGroup10: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_361_store_0_req_0;
      ptr_deref_361_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_361_store_0_req_1;
      ptr_deref_361_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup10_gI: SplitGuardInterface generic map(name => "StoreGroup10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_361_word_address_0;
      data_in <= ptr_deref_361_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup10 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_14_sr_req(0),
          mack => memory_space_14_sr_ack(0),
          maddr => memory_space_14_sr_addr(0 downto 0),
          mdata => memory_space_14_sr_data(31 downto 0),
          mtag => memory_space_14_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup10 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_14_sc_req(0),
          mack => memory_space_14_sc_ack(0),
          mtag => memory_space_14_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 10
    -- shared store operator group (11) : ptr_deref_78_store_0 
    StoreGroup11: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_78_store_0_req_0;
      ptr_deref_78_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_78_store_0_req_1;
      ptr_deref_78_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup11_gI: SplitGuardInterface generic map(name => "StoreGroup11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_78_word_address_0;
      data_in <= ptr_deref_78_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup11 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(0 downto 0),
          mdata => memory_space_9_sr_data(15 downto 0),
          mtag => memory_space_9_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup11 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 11
    -- shared store operator group (12) : ptr_deref_92_store_0 
    StoreGroup12: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_92_store_0_req_0;
      ptr_deref_92_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_92_store_0_req_1;
      ptr_deref_92_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup12_gI: SplitGuardInterface generic map(name => "StoreGroup12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_92_word_address_0;
      data_in <= ptr_deref_92_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup12 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(0 downto 0),
          mdata => memory_space_10_sr_data(31 downto 0),
          mtag => memory_space_10_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup12 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 12
    -- shared inport operator group (0) : RPIPE_ebbyNo_in_89_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_ebbyNo_in_89_inst_req_0;
      RPIPE_ebbyNo_in_89_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_ebbyNo_in_89_inst_req_1;
      RPIPE_ebbyNo_in_89_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_6_90 <= data_out(31 downto 0);
      ebbyNo_in_read_0_gI: SplitGuardInterface generic map(name => "ebbyNo_in_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ebbyNo_in_read_0: InputPortRevised -- 
        generic map ( name => "ebbyNo_in_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ebbyNo_in_pipe_read_req(0),
          oack => ebbyNo_in_pipe_read_ack(0),
          odata => ebbyNo_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_matrix_in_300_inst RPIPE_matrix_in_136_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_matrix_in_300_inst_req_0;
      reqL_unguarded(0) <= RPIPE_matrix_in_136_inst_req_0;
      RPIPE_matrix_in_300_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_matrix_in_136_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_matrix_in_300_inst_req_1;
      reqR_unguarded(0) <= RPIPE_matrix_in_136_inst_req_1;
      RPIPE_matrix_in_300_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_matrix_in_136_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      iNsTr_57_301 <= data_out(31 downto 16);
      iNsTr_17_137 <= data_out(15 downto 0);
      matrix_in_read_1_gI: SplitGuardInterface generic map(name => "matrix_in_read_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      matrix_in_read_1: InputPortRevised -- 
        generic map ( name => "matrix_in_read_1", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => matrix_in_pipe_read_req(0),
          oack => matrix_in_pipe_read_ack(0),
          odata => matrix_in_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_maxNitr_in_75_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_maxNitr_in_75_inst_req_0;
      RPIPE_maxNitr_in_75_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_maxNitr_in_75_inst_req_1;
      RPIPE_maxNitr_in_75_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_1_76 <= data_out(15 downto 0);
      maxNitr_in_read_2_gI: SplitGuardInterface generic map(name => "maxNitr_in_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxNitr_in_read_2: InputPortRevised -- 
        generic map ( name => "maxNitr_in_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxNitr_in_pipe_read_req(0),
          oack => maxNitr_in_pipe_read_ack(0),
          odata => maxNitr_in_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_rate_in_358_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_rate_in_358_inst_req_0;
      RPIPE_rate_in_358_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_rate_in_358_inst_req_1;
      RPIPE_rate_in_358_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_68_359 <= data_out(31 downto 0);
      rate_in_read_3_gI: SplitGuardInterface generic map(name => "rate_in_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      rate_in_read_3: InputPortRevised -- 
        generic map ( name => "rate_in_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => rate_in_pipe_read_req(0),
          oack => rate_in_pipe_read_ack(0),
          odata => rate_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_10: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_10",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_10_lr_addr,
      lr_req_in => memory_space_10_lr_req,
      lr_ack_out => memory_space_10_lr_ack,
      lr_tag_in => memory_space_10_lr_tag,
      lc_req_in => memory_space_10_lc_req,
      lc_ack_out => memory_space_10_lc_ack,
      lc_data_out => memory_space_10_lc_data,
      lc_tag_out => memory_space_10_lc_tag,
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_11: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_11",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_11_lr_addr,
      lr_req_in => memory_space_11_lr_req,
      lr_ack_out => memory_space_11_lr_ack,
      lr_tag_in => memory_space_11_lr_tag,
      lc_req_in => memory_space_11_lc_req,
      lc_ack_out => memory_space_11_lc_ack,
      lc_data_out => memory_space_11_lc_data,
      lc_tag_out => memory_space_11_lc_tag,
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_12: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_12",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_12_lr_addr,
      lr_req_in => memory_space_12_lr_req,
      lr_ack_out => memory_space_12_lr_ack,
      lr_tag_in => memory_space_12_lr_tag,
      lc_req_in => memory_space_12_lc_req,
      lc_ack_out => memory_space_12_lc_ack,
      lc_data_out => memory_space_12_lc_data,
      lc_tag_out => memory_space_12_lc_tag,
      sr_addr_in => memory_space_12_sr_addr,
      sr_data_in => memory_space_12_sr_data,
      sr_req_in => memory_space_12_sr_req,
      sr_ack_out => memory_space_12_sr_ack,
      sr_tag_in => memory_space_12_sr_tag,
      sc_req_in=> memory_space_12_sc_req,
      sc_ack_out => memory_space_12_sc_ack,
      sc_tag_out => memory_space_12_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_13: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_13",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_13_lr_addr,
      lr_req_in => memory_space_13_lr_req,
      lr_ack_out => memory_space_13_lr_ack,
      lr_tag_in => memory_space_13_lr_tag,
      lc_req_in => memory_space_13_lc_req,
      lc_ack_out => memory_space_13_lc_ack,
      lc_data_out => memory_space_13_lc_data,
      lc_tag_out => memory_space_13_lc_tag,
      sr_addr_in => memory_space_13_sr_addr,
      sr_data_in => memory_space_13_sr_data,
      sr_req_in => memory_space_13_sr_req,
      sr_ack_out => memory_space_13_sr_ack,
      sr_tag_in => memory_space_13_sr_tag,
      sc_req_in=> memory_space_13_sc_req,
      sc_ack_out => memory_space_13_sc_ack,
      sc_tag_out => memory_space_13_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_14: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_14",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_14_lr_addr,
      lr_req_in => memory_space_14_lr_req,
      lr_ack_out => memory_space_14_lr_ack,
      lr_tag_in => memory_space_14_lr_tag,
      lc_req_in => memory_space_14_lc_req,
      lc_ack_out => memory_space_14_lc_ack,
      lc_data_out => memory_space_14_lc_data,
      lc_tag_out => memory_space_14_lc_tag,
      sr_addr_in => memory_space_14_sr_addr,
      sr_data_in => memory_space_14_sr_data,
      sr_req_in => memory_space_14_sr_req,
      sr_ack_out => memory_space_14_sr_ack,
      sr_tag_in => memory_space_14_sr_tag,
      sc_req_in=> memory_space_14_sc_req,
      sc_ack_out => memory_space_14_sc_ack,
      sc_tag_out => memory_space_14_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_9",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end initInputs_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity initialize_aPriori is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initialize_aPriori;
architecture initialize_aPriori_arch of initialize_aPriori is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal initialize_aPriori_CP_2378_start: Boolean;
  signal initialize_aPriori_CP_2378_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_402_inst_req_0 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal ptr_deref_383_store_0_ack_0 : boolean;
  signal LOAD_ncols_398_load_0_ack_0 : boolean;
  signal ptr_deref_383_store_0_req_0 : boolean;
  signal LOAD_ncols_398_load_0_req_0 : boolean;
  signal SLT_i32_u1_409_inst_ack_0 : boolean;
  signal type_cast_402_inst_ack_1 : boolean;
  signal LOAD_ncols_398_load_0_ack_1 : boolean;
  signal LOAD_ncols_398_load_0_req_1 : boolean;
  signal type_cast_402_inst_req_1 : boolean;
  signal ptr_deref_391_load_0_ack_1 : boolean;
  signal type_cast_402_inst_ack_0 : boolean;
  signal SLT_i32_u1_409_inst_req_0 : boolean;
  signal ptr_deref_420_load_0_req_1 : boolean;
  signal ptr_deref_420_load_0_ack_0 : boolean;
  signal ptr_deref_383_store_0_req_1 : boolean;
  signal ptr_deref_383_store_0_ack_1 : boolean;
  signal ptr_deref_391_load_0_req_0 : boolean;
  signal if_stmt_411_branch_ack_0 : boolean;
  signal ptr_deref_391_load_0_ack_0 : boolean;
  signal SLT_i32_u1_409_inst_req_1 : boolean;
  signal if_stmt_411_branch_req_0 : boolean;
  signal SLT_i32_u1_409_inst_ack_1 : boolean;
  signal ptr_deref_420_load_0_ack_1 : boolean;
  signal type_cast_424_inst_req_0 : boolean;
  signal type_cast_424_inst_ack_0 : boolean;
  signal ptr_deref_420_load_0_req_0 : boolean;
  signal ptr_deref_391_load_0_req_1 : boolean;
  signal ptr_deref_428_load_0_req_0 : boolean;
  signal type_cast_424_inst_req_1 : boolean;
  signal type_cast_424_inst_ack_1 : boolean;
  signal type_cast_432_inst_req_0 : boolean;
  signal type_cast_432_inst_ack_0 : boolean;
  signal type_cast_432_inst_req_1 : boolean;
  signal type_cast_432_inst_ack_1 : boolean;
  signal if_stmt_411_branch_ack_1 : boolean;
  signal ptr_deref_428_load_0_ack_0 : boolean;
  signal ptr_deref_428_load_0_req_1 : boolean;
  signal ptr_deref_428_load_0_ack_1 : boolean;
  signal addr_of_437_final_reg_req_0 : boolean;
  signal addr_of_437_final_reg_ack_0 : boolean;
  signal addr_of_437_final_reg_req_1 : boolean;
  signal addr_of_437_final_reg_ack_1 : boolean;
  signal ptr_deref_440_store_0_req_0 : boolean;
  signal ptr_deref_440_store_0_ack_0 : boolean;
  signal ptr_deref_440_store_0_req_1 : boolean;
  signal ptr_deref_440_store_0_ack_1 : boolean;
  signal ptr_deref_447_load_0_req_0 : boolean;
  signal ptr_deref_447_load_0_ack_0 : boolean;
  signal ptr_deref_447_load_0_req_1 : boolean;
  signal ptr_deref_447_load_0_ack_1 : boolean;
  signal ADD_u16_u16_453_inst_req_0 : boolean;
  signal ADD_u16_u16_453_inst_ack_0 : boolean;
  signal ADD_u16_u16_453_inst_req_1 : boolean;
  signal ADD_u16_u16_453_inst_ack_1 : boolean;
  signal ptr_deref_456_store_0_req_0 : boolean;
  signal ptr_deref_456_store_0_ack_0 : boolean;
  signal ptr_deref_456_store_0_req_1 : boolean;
  signal ptr_deref_456_store_0_ack_1 : boolean;
  signal memory_space_15_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_15_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_15_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_15_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_15_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_15_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_15_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_sc_tag :  std_logic_vector(2 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initialize_aPriori_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initialize_aPriori_CP_2378_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initialize_aPriori_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initialize_aPriori_CP_2378_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initialize_aPriori_CP_2378_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initialize_aPriori_CP_2378_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initialize_aPriori_CP_2378: Block -- control-path 
    signal initialize_aPriori_CP_2378_elements: BooleanArray(75 downto 0);
    -- 
  begin -- 
    initialize_aPriori_CP_2378_elements(0) <= initialize_aPriori_CP_2378_start;
    initialize_aPriori_CP_2378_symbol <= initialize_aPriori_CP_2378_elements(75);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_376/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_376/branch_block_stmt_376__entry__
      -- CP-element group 1: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386__entry__
      -- 
    initialize_aPriori_CP_2378_elements(1) <= initialize_aPriori_CP_2378_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386__exit__
      -- CP-element group 2: 	 branch_block_stmt_376/bb_0_bb_1
      -- 
    initialize_aPriori_CP_2378_elements(2) <= initialize_aPriori_CP_2378_elements(13);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	62 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	14 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410__entry__
      -- CP-element group 3: 	 branch_block_stmt_376/merge_stmt_388__exit__
      -- 
    initialize_aPriori_CP_2378_elements(3) <= initialize_aPriori_CP_2378_elements(62);
    -- CP-element group 4:  branch  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	25 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	26 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_376/if_stmt_411__entry__
      -- CP-element group 4: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410__exit__
      -- 
    initialize_aPriori_CP_2378_elements(4) <= initialize_aPriori_CP_2378_elements(25);
    -- CP-element group 5:  merge  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	65 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	35 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442__entry__
      -- CP-element group 5: 	 branch_block_stmt_376/merge_stmt_417__exit__
      -- 
    initialize_aPriori_CP_2378_elements(5) <= initialize_aPriori_CP_2378_elements(65);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	49 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	66 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_376/bb_2_bb_3
      -- CP-element group 6: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442__exit__
      -- 
    initialize_aPriori_CP_2378_elements(6) <= initialize_aPriori_CP_2378_elements(49);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	68 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	50 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458__entry__
      -- CP-element group 7: 	 branch_block_stmt_376/merge_stmt_444__exit__
      -- 
    initialize_aPriori_CP_2378_elements(7) <= initialize_aPriori_CP_2378_elements(68);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	57 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	60 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_376/bb_3_bb_1
      -- CP-element group 8: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458__exit__
      -- 
    initialize_aPriori_CP_2378_elements(8) <= initialize_aPriori_CP_2378_elements(57);
    -- CP-element group 9:  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	71 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	72 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_376/return__
      -- CP-element group 9: 	 branch_block_stmt_376/merge_stmt_460__exit__
      -- 
    initialize_aPriori_CP_2378_elements(9) <= initialize_aPriori_CP_2378_elements(71);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	74 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	75 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_376/branch_block_stmt_376__exit__
      -- CP-element group 10: 	 branch_block_stmt_376/merge_stmt_462__exit__
      -- 
    initialize_aPriori_CP_2378_elements(10) <= initialize_aPriori_CP_2378_elements(74);
    -- CP-element group 11:  fork  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (31) 
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_word_addrgen/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/word_0/rr
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_word_addrgen/$exit
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_addr_resize/base_resize_ack
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_word_addrgen/root_register_req
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_addr_resize/base_resize_req
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_word_addrgen/root_register_ack
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_addr_resize/$exit
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_addr_resize/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/word_0/cr
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/word_0/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_base_address_resized
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/ptr_deref_383_Split/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/ptr_deref_383_Split/$exit
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_update_start_
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/ptr_deref_383_Split/split_req
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/ptr_deref_383_Split/split_ack
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/$entry
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_root_address_calculated
      -- 
    cr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(11), ack => ptr_deref_383_store_0_req_1); -- 
    rr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(11), ack => ptr_deref_383_store_0_req_0); -- 
    initialize_aPriori_CP_2378_elements(11) <= initialize_aPriori_CP_2378_elements(1);
    -- CP-element group 12:  transition  input  no-bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/word_0/ra
      -- CP-element group 12: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_sample_completed_
      -- 
    ra_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_store_0_ack_0, ack => initialize_aPriori_CP_2378_elements(12)); -- 
    -- CP-element group 13:  transition  input  no-bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	2 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/$exit
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_376/assign_stmt_381_to_assign_stmt_386/ptr_deref_383_update_completed_
      -- 
    ca_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_383_store_0_ack_1, ack => initialize_aPriori_CP_2378_elements(13)); -- 
    -- CP-element group 14:  join  fork  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	3 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	22 
    -- CP-element group 14: 	25 
    -- CP-element group 14:  members (48) 
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_update_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_update_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_root_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_update_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_word_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/word_0/cr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_update_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_update_start_
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_word_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_root_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_address_resized
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_addr_resize/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_addr_resize/$exit
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_plus_offset/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_plus_offset/$exit
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_word_addrgen/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_word_addrgen/$exit
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_word_addrgen/root_register_req
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/word_0/cr
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_word_addrgen/root_register_ack
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_sample_start_
      -- 
    cr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => ptr_deref_391_load_0_req_1); -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => ptr_deref_391_load_0_req_0); -- 
    cr_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => type_cast_395_inst_req_1); -- 
    cr_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => LOAD_ncols_398_load_0_req_1); -- 
    rr_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => LOAD_ncols_398_load_0_req_0); -- 
    cr_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => type_cast_402_inst_req_1); -- 
    cr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(14), ack => SLT_i32_u1_409_inst_req_1); -- 
    initialize_aPriori_CP_2378_elements(14) <= initialize_aPriori_CP_2378_elements(3);
    -- CP-element group 15:  transition  input  no-bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Sample/word_access_start/word_0/ra
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_391_load_0_ack_0, ack => initialize_aPriori_CP_2378_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  no-bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/ptr_deref_391_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/ptr_deref_391_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/ptr_deref_391_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/ptr_deref_391_Update/ptr_deref_391_Merge/$entry
      -- 
    ca_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_391_load_0_ack_1, ack => initialize_aPriori_CP_2378_elements(16)); -- 
    rr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(16), ack => type_cast_395_inst_req_0); -- 
    -- CP-element group 17:  transition  input  no-bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Sample/ra
      -- 
    ra_2520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(17)); -- 
    -- CP-element group 18:  transition  input  no-bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_395_Update/$exit
      -- 
    ca_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(18)); -- 
    -- CP-element group 19:  transition  input  no-bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	14 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_sample_completed_
      -- 
    ra_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_398_load_0_ack_0, ack => initialize_aPriori_CP_2378_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  no-bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/LOAD_ncols_398_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/LOAD_ncols_398_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/LOAD_ncols_398_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/LOAD_ncols_398_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/LOAD_ncols_398_Update/word_access_complete/$exit
      -- 
    ca_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_398_load_0_ack_1, ack => initialize_aPriori_CP_2378_elements(20)); -- 
    rr_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(20), ack => type_cast_402_inst_req_0); -- 
    -- CP-element group 21:  transition  input  no-bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Sample/ra
      -- 
    ra_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(21)); -- 
    -- CP-element group 22:  transition  input  no-bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	14 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/type_cast_402_Update/ca
      -- 
    ca_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Sample/rr
      -- 
    rr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(23), ack => SLT_i32_u1_409_inst_req_0); -- 
    initialize_aPriori_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "initialize_aPriori_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialize_aPriori_CP_2378_elements(18) & initialize_aPriori_CP_2378_elements(22);
      gj_initialize_aPriori_cp_element_group_23 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialize_aPriori_CP_2378_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  no-bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Sample/ra
      -- 
    ra_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_409_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(24)); -- 
    -- CP-element group 25:  transition  input  no-bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	14 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	4 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/$exit
      -- CP-element group 25: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_376/assign_stmt_392_to_assign_stmt_410/SLT_i32_u1_409_Update/ca
      -- 
    ca_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_409_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(25)); -- 
    -- CP-element group 26:  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	4 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_376/if_stmt_411_dead_link/$entry
      -- 
    initialize_aPriori_CP_2378_elements(26) <= initialize_aPriori_CP_2378_elements(4);
    -- CP-element group 27:  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_376/if_stmt_411_eval_test/branch_req
      -- CP-element group 27: 	 branch_block_stmt_376/if_stmt_411_eval_test/$entry
      -- CP-element group 27: 	 branch_block_stmt_376/if_stmt_411_eval_test/$exit
      -- 
    branch_req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(27), ack => if_stmt_411_branch_req_0); -- 
    initialize_aPriori_CP_2378_elements(27) <= initialize_aPriori_CP_2378_elements(4);
    -- CP-element group 28:  branch  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_376/R_iNsTr_6_412_place
      -- 
    initialize_aPriori_CP_2378_elements(28) <= initialize_aPriori_CP_2378_elements(27);
    -- CP-element group 29:  transition  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_376/if_stmt_411_if_link/$entry
      -- 
    initialize_aPriori_CP_2378_elements(29) <= initialize_aPriori_CP_2378_elements(28);
    -- CP-element group 30:  transition  input  no-bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_376/if_stmt_411_if_link/if_choice_transition
      -- CP-element group 30: 	 branch_block_stmt_376/if_stmt_411_if_link/$exit
      -- 
    if_choice_transition_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_411_branch_ack_1, ack => initialize_aPriori_CP_2378_elements(30)); -- 
    -- CP-element group 31:  transition  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	28 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_376/if_stmt_411_else_link/$entry
      -- 
    initialize_aPriori_CP_2378_elements(31) <= initialize_aPriori_CP_2378_elements(28);
    -- CP-element group 32:  transition  input  no-bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_376/if_stmt_411_else_link/else_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_376/if_stmt_411_else_link/$exit
      -- 
    else_choice_transition_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_411_branch_ack_0, ack => initialize_aPriori_CP_2378_elements(32)); -- 
    -- CP-element group 33:  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	63 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_376/bb_1_bb_2
      -- 
    initialize_aPriori_CP_2378_elements(33) <= initialize_aPriori_CP_2378_elements(30);
    -- CP-element group 34:  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	69 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_376/bb_1_bb_4
      -- 
    initialize_aPriori_CP_2378_elements(34) <= initialize_aPriori_CP_2378_elements(32);
    -- CP-element group 35:  join  fork  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	5 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	39 
    -- CP-element group 35: 	40 
    -- CP-element group 35: 	41 
    -- CP-element group 35: 	43 
    -- CP-element group 35: 	45 
    -- CP-element group 35: 	48 
    -- CP-element group 35:  members (67) 
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/word_0/cr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_word_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_address_resized
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_word_addrgen/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_word_addrgen/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_addr_resize/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_base_addr_resize/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_word_addrgen/root_register_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/word_0/rr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_word_addrgen/root_register_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_addr_resize/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_addr_resize/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/word_0/rr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_word_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_address_resized
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/word_0/cr
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_word_addrgen/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_word_addrgen/$exit
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_word_addrgen/root_register_req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_word_addrgen/root_register_ack
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_complete/req
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_update_start_
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/word_0/cr
      -- 
    cr_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => ptr_deref_420_load_0_req_1); -- 
    rr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => ptr_deref_420_load_0_req_0); -- 
    cr_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => type_cast_424_inst_req_1); -- 
    cr_2716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => ptr_deref_428_load_0_req_1); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => ptr_deref_428_load_0_req_0); -- 
    cr_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => type_cast_432_inst_req_1); -- 
    req_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => addr_of_437_final_reg_req_1); -- 
    cr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(35), ack => ptr_deref_440_store_0_req_1); -- 
    initialize_aPriori_CP_2378_elements(35) <= initialize_aPriori_CP_2378_elements(5);
    -- CP-element group 36:  transition  input  no-bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/word_0/ra
      -- CP-element group 36: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Sample/$exit
      -- 
    ra_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_420_load_0_ack_0, ack => initialize_aPriori_CP_2378_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  no-bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (12) 
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/ptr_deref_420_Merge/merge_ack
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/ptr_deref_420_Merge/merge_req
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/ptr_deref_420_Merge/$entry
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/ptr_deref_420_Merge/$exit
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_420_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_sample_start_
      -- 
    ca_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_420_load_0_ack_1, ack => initialize_aPriori_CP_2378_elements(37)); -- 
    rr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(37), ack => type_cast_424_inst_req_0); -- 
    -- CP-element group 38:  transition  input  no-bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_sample_completed_
      -- 
    ra_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(38)); -- 
    -- CP-element group 39:  transition  input  no-bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	35 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	46 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_424_Update/ca
      -- 
    ca_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(39)); -- 
    -- CP-element group 40:  transition  input  no-bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Sample/word_access_start/word_0/ra
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_428_load_0_ack_0, ack => initialize_aPriori_CP_2378_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  no-bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	35 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (12) 
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/ptr_deref_428_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/ptr_deref_428_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/ptr_deref_428_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_428_Update/ptr_deref_428_Merge/merge_ack
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Sample/$entry
      -- 
    ca_2717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_428_load_0_ack_1, ack => initialize_aPriori_CP_2378_elements(41)); -- 
    rr_2730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(41), ack => type_cast_432_inst_req_0); -- 
    -- CP-element group 42:  transition  input  no-bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Sample/$exit
      -- 
    ra_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  no-bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	35 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (27) 
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_scaled_0
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_computed_0
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_resize_0/$entry
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_resize_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_resize_0/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_resize_0/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_scale_0/$entry
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_scale_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_scale_0/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_scale_0/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_final_index_sum_regn/$entry
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_final_index_sum_regn/$exit
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_offset_calculated
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_index_resized_0
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/type_cast_432_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_final_index_sum_regn/req
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_final_index_sum_regn/ack
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/array_obj_ref_436_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_request/$entry
      -- CP-element group 43: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_request/req
      -- 
    ca_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(43)); -- 
    req_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(43), ack => addr_of_437_final_reg_req_0); -- 
    -- CP-element group 44:  transition  input  no-bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	49 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_request/$exit
      -- CP-element group 44: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_request/ack
      -- 
    ack_2770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_437_final_reg_ack_0, ack => initialize_aPriori_CP_2378_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  no-bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	35 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (19) 
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/addr_of_437_complete/ack
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_word_addrgen/root_register_ack
      -- 
    ack_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_437_final_reg_ack_1, ack => initialize_aPriori_CP_2378_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	39 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/ptr_deref_440_Split/$entry
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/ptr_deref_440_Split/$exit
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/ptr_deref_440_Split/split_req
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/ptr_deref_440_Split/split_ack
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/word_0/rr
      -- 
    rr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(46), ack => ptr_deref_440_store_0_req_0); -- 
    initialize_aPriori_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "initialize_aPriori_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialize_aPriori_CP_2378_elements(39) & initialize_aPriori_CP_2378_elements(45);
      gj_initialize_aPriori_cp_element_group_46 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialize_aPriori_CP_2378_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  no-bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Sample/word_access_start/word_0/ra
      -- 
    ra_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_440_store_0_ack_0, ack => initialize_aPriori_CP_2378_elements(47)); -- 
    -- CP-element group 48:  transition  input  no-bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/ptr_deref_440_Update/word_access_complete/word_0/ca
      -- 
    ca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_440_store_0_ack_1, ack => initialize_aPriori_CP_2378_elements(48)); -- 
    -- CP-element group 49:  join  transition  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	44 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	6 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_376/assign_stmt_421_to_assign_stmt_442/$exit
      -- 
    initialize_aPriori_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "initialize_aPriori_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initialize_aPriori_CP_2378_elements(44) & initialize_aPriori_CP_2378_elements(48);
      gj_initialize_aPriori_cp_element_group_49 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialize_aPriori_CP_2378_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  fork  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	7 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	55 
    -- CP-element group 50: 	57 
    -- CP-element group 50:  members (51) 
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_update_start_
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_word_addrgen/root_register_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/word_0/rr
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/word_0/cr
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_update_start_
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Update/cr
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_update_start_
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_word_addrgen/root_register_ack
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/word_0/cr
      -- 
    cr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(50), ack => ptr_deref_447_load_0_req_1); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(50), ack => ptr_deref_447_load_0_req_0); -- 
    cr_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(50), ack => ADD_u16_u16_453_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(50), ack => ptr_deref_456_store_0_req_1); -- 
    initialize_aPriori_CP_2378_elements(50) <= initialize_aPriori_CP_2378_elements(7);
    -- CP-element group 51:  transition  input  no-bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	58 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Sample/word_access_start/word_0/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_447_load_0_ack_0, ack => initialize_aPriori_CP_2378_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  no-bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/word_access_complete/word_0/ca
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/ptr_deref_447_Merge/$entry
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/ptr_deref_447_Merge/$exit
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/ptr_deref_447_Merge/merge_req
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_Update/ptr_deref_447_Merge/merge_ack
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Sample/rr
      -- 
    ca_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_447_load_0_ack_1, ack => initialize_aPriori_CP_2378_elements(52)); -- 
    rr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(52), ack => ADD_u16_u16_453_inst_req_0); -- 
    -- CP-element group 53:  transition  input  no-bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Sample/ra
      -- 
    ra_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_453_inst_ack_0, ack => initialize_aPriori_CP_2378_elements(53)); -- 
    -- CP-element group 54:  transition  input  no-bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	50 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ADD_u16_u16_453_Update/ca
      -- 
    ca_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_453_inst_ack_1, ack => initialize_aPriori_CP_2378_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  no-bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	58 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/ptr_deref_456_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/ptr_deref_456_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/ptr_deref_456_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/ptr_deref_456_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/word_0/rr
      -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initialize_aPriori_CP_2378_elements(55), ack => ptr_deref_456_store_0_req_0); -- 
    initialize_aPriori_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 38) := "initialize_aPriori_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initialize_aPriori_CP_2378_elements(50) & initialize_aPriori_CP_2378_elements(54) & initialize_aPriori_CP_2378_elements(58);
      gj_initialize_aPriori_cp_element_group_55 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initialize_aPriori_CP_2378_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  no-bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Sample/word_access_start/word_0/ra
      -- 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_456_store_0_ack_0, ack => initialize_aPriori_CP_2378_elements(56)); -- 
    -- CP-element group 57:  transition  input  no-bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	50 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	8 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/$exit
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_456_Update/word_access_complete/word_0/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_456_store_0_ack_1, ack => initialize_aPriori_CP_2378_elements(57)); -- 
    -- CP-element group 58:  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	55 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_376/assign_stmt_448_to_assign_stmt_458/ptr_deref_447_ptr_deref_456_delay
      -- 
    -- Element group initialize_aPriori_CP_2378_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => initialize_aPriori_CP_2378_elements(51), ack => initialize_aPriori_CP_2378_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  transition  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_376/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_376/bb_0_bb_1_PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(59) <= initialize_aPriori_CP_2378_elements(2);
    -- CP-element group 60:  transition  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	8 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_376/bb_3_bb_1_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_376/bb_3_bb_1_PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(60) <= initialize_aPriori_CP_2378_elements(8);
    -- CP-element group 61:  merge  place  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_376/merge_stmt_388_PhiReqMerge
      -- 
    initialize_aPriori_CP_2378_elements(61) <= OrReduce(initialize_aPriori_CP_2378_elements(59) & initialize_aPriori_CP_2378_elements(60));
    -- CP-element group 62:  transition  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	3 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_376/merge_stmt_388_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_376/merge_stmt_388_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_376/merge_stmt_388_PhiAck/dummy
      -- 
    initialize_aPriori_CP_2378_elements(62) <= initialize_aPriori_CP_2378_elements(61);
    -- CP-element group 63:  transition  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	33 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_376/bb_1_bb_2_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_376/bb_1_bb_2_PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(63) <= initialize_aPriori_CP_2378_elements(33);
    -- CP-element group 64:  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_376/merge_stmt_417_PhiReqMerge
      -- 
    initialize_aPriori_CP_2378_elements(64) <= initialize_aPriori_CP_2378_elements(63);
    -- CP-element group 65:  transition  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	5 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_376/merge_stmt_417_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_376/merge_stmt_417_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_376/merge_stmt_417_PhiAck/dummy
      -- 
    initialize_aPriori_CP_2378_elements(65) <= initialize_aPriori_CP_2378_elements(64);
    -- CP-element group 66:  transition  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	6 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_376/bb_2_bb_3_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_376/bb_2_bb_3_PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(66) <= initialize_aPriori_CP_2378_elements(6);
    -- CP-element group 67:  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_376/merge_stmt_444_PhiReqMerge
      -- 
    initialize_aPriori_CP_2378_elements(67) <= initialize_aPriori_CP_2378_elements(66);
    -- CP-element group 68:  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	7 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_376/merge_stmt_444_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_376/merge_stmt_444_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_376/merge_stmt_444_PhiAck/dummy
      -- 
    initialize_aPriori_CP_2378_elements(68) <= initialize_aPriori_CP_2378_elements(67);
    -- CP-element group 69:  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	34 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_376/bb_1_bb_4_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_376/bb_1_bb_4_PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(69) <= initialize_aPriori_CP_2378_elements(34);
    -- CP-element group 70:  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_376/merge_stmt_460_PhiReqMerge
      -- 
    initialize_aPriori_CP_2378_elements(70) <= initialize_aPriori_CP_2378_elements(69);
    -- CP-element group 71:  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	9 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_376/merge_stmt_460_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_376/merge_stmt_460_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_376/merge_stmt_460_PhiAck/dummy
      -- 
    initialize_aPriori_CP_2378_elements(71) <= initialize_aPriori_CP_2378_elements(70);
    -- CP-element group 72:  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_376/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_376/return___PhiReq/$exit
      -- 
    initialize_aPriori_CP_2378_elements(72) <= initialize_aPriori_CP_2378_elements(9);
    -- CP-element group 73:  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_376/merge_stmt_462_PhiReqMerge
      -- 
    initialize_aPriori_CP_2378_elements(73) <= initialize_aPriori_CP_2378_elements(72);
    -- CP-element group 74:  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	10 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_376/merge_stmt_462_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_376/merge_stmt_462_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_376/merge_stmt_462_PhiAck/dummy
      -- 
    initialize_aPriori_CP_2378_elements(74) <= initialize_aPriori_CP_2378_elements(73);
    -- CP-element group 75:  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	10 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_376/$exit
      -- CP-element group 75: 	 $exit
      -- 
    initialize_aPriori_CP_2378_elements(75) <= initialize_aPriori_CP_2378_elements(10);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_381 : std_logic_vector(31 downto 0);
    signal LOAD_ncols_398_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_398_word_address_0 : std_logic_vector(0 downto 0);
    signal R_iNsTr_12_435_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_12_435_scaled : std_logic_vector(9 downto 0);
    signal array_obj_ref_436_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_436_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_436_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_436_root_address : std_logic_vector(9 downto 0);
    signal iNsTr_10_425 : std_logic_vector(31 downto 0);
    signal iNsTr_11_429 : std_logic_vector(15 downto 0);
    signal iNsTr_12_433 : std_logic_vector(63 downto 0);
    signal iNsTr_13_438 : std_logic_vector(31 downto 0);
    signal iNsTr_17_448 : std_logic_vector(15 downto 0);
    signal iNsTr_18_454 : std_logic_vector(15 downto 0);
    signal iNsTr_2_392 : std_logic_vector(15 downto 0);
    signal iNsTr_3_396 : std_logic_vector(31 downto 0);
    signal iNsTr_4_399 : std_logic_vector(15 downto 0);
    signal iNsTr_5_403 : std_logic_vector(31 downto 0);
    signal iNsTr_6_410 : std_logic_vector(0 downto 0);
    signal iNsTr_9_421 : std_logic_vector(15 downto 0);
    signal ptr_deref_383_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_383_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_383_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_383_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_383_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_383_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_391_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_391_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_391_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_391_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_391_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_420_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_420_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_420_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_420_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_420_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_428_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_428_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_428_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_428_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_428_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_440_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_440_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_440_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_440_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_440_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_440_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_447_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_447_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_447_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_447_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_447_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_456_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_456_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_456_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_456_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_456_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_456_word_offset_0 : std_logic_vector(0 downto 0);
    signal type_cast_385_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_406_wire : std_logic_vector(31 downto 0);
    signal type_cast_408_wire : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(15 downto 0);
    signal xxinitialize_aPriorixxbodyxxI_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    I_381 <= "00000000000000000000000000000000";
    LOAD_ncols_398_word_address_0 <= "0";
    array_obj_ref_436_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_436_resized_base_address <= "0000000000";
    ptr_deref_383_word_offset_0 <= "0";
    ptr_deref_391_word_offset_0 <= "0";
    ptr_deref_420_word_offset_0 <= "0";
    ptr_deref_428_word_offset_0 <= "0";
    ptr_deref_440_word_offset_0 <= "0000000000";
    ptr_deref_447_word_offset_0 <= "0";
    ptr_deref_456_word_offset_0 <= "0";
    type_cast_385_wire_constant <= "0000000000000000";
    type_cast_452_wire_constant <= "0000000000000001";
    xxinitialize_aPriorixxbodyxxI_alloc_base_address <= "0";
    addr_of_437_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_437_final_reg_req_0;
      addr_of_437_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_437_final_reg_req_1;
      addr_of_437_final_reg_ack_1<= rack(0);
      addr_of_437_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_437_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_436_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_13_438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_2_392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_3_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_402_inst_req_0;
      type_cast_402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_402_inst_req_1;
      type_cast_402_inst_ack_1<= rack(0);
      type_cast_402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_4_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_5_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_406_inst
    process(iNsTr_3_396) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_3_396(31 downto 0);
      type_cast_406_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_408_inst
    process(iNsTr_5_403) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_5_403(31 downto 0);
      type_cast_408_wire <= tmp_var; -- 
    end process;
    type_cast_432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_432_inst_req_0;
      type_cast_432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_432_inst_req_1;
      type_cast_432_inst_ack_1<= rack(0);
      type_cast_432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_11_429,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_12_433,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_ncols_398_gather_scatter
    process(LOAD_ncols_398_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_398_data_0;
      ov(15 downto 0) := iv;
      iNsTr_4_399 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_436_index_0_rename
    process(R_iNsTr_12_435_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_12_435_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_12_435_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_436_index_0_resize
    process(iNsTr_12_433) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_12_433;
      ov := iv(9 downto 0);
      R_iNsTr_12_435_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_436_index_offset
    process(R_iNsTr_12_435_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_12_435_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_436_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_436_root_address_inst
    process(array_obj_ref_436_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_436_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_436_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_addr_0
    process(ptr_deref_383_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_383_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_383_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_gather_scatter
    process(type_cast_385_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_385_wire_constant;
      ov(15 downto 0) := iv;
      ptr_deref_383_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_383_root_address_inst
    process(ptr_deref_383_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_383_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_383_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_391_addr_0
    process(ptr_deref_391_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_391_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_391_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_391_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_391_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_391_gather_scatter
    process(ptr_deref_391_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_391_data_0;
      ov(15 downto 0) := iv;
      iNsTr_2_392 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_391_root_address_inst
    process(ptr_deref_391_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_391_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_391_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_addr_0
    process(ptr_deref_420_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_420_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_420_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_420_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_gather_scatter
    process(ptr_deref_420_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_420_data_0;
      ov(15 downto 0) := iv;
      iNsTr_9_421 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_root_address_inst
    process(ptr_deref_420_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_420_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_420_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_428_addr_0
    process(ptr_deref_428_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_428_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_428_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_428_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_428_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_428_gather_scatter
    process(ptr_deref_428_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_428_data_0;
      ov(15 downto 0) := iv;
      iNsTr_11_429 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_428_root_address_inst
    process(ptr_deref_428_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_428_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_428_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_440_addr_0
    process(ptr_deref_440_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_440_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_440_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_440_base_resize
    process(iNsTr_13_438) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_438;
      ov := iv(9 downto 0);
      ptr_deref_440_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_440_gather_scatter
    process(iNsTr_10_425) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_425;
      ov(31 downto 0) := iv;
      ptr_deref_440_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_440_root_address_inst
    process(ptr_deref_440_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_440_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_440_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_addr_0
    process(ptr_deref_447_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_447_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_447_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_gather_scatter
    process(ptr_deref_447_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_data_0;
      ov(15 downto 0) := iv;
      iNsTr_17_448 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_root_address_inst
    process(ptr_deref_447_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_447_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_addr_0
    process(ptr_deref_456_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_456_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_456_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_base_resize
    process(I_381) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_381;
      ov := iv(0 downto 0);
      ptr_deref_456_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_gather_scatter
    process(iNsTr_18_454) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_454;
      ov(15 downto 0) := iv;
      ptr_deref_456_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_root_address_inst
    process(ptr_deref_456_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_456_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_456_root_address <= ov(0 downto 0);
      --
    end process;
    if_stmt_411_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_6_410;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_411_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_411_branch_req_0,
          ack0 => if_stmt_411_branch_ack_0,
          ack1 => if_stmt_411_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u16_u16_453_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_17_448;
      iNsTr_18_454 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_453_inst_req_0;
      ADD_u16_u16_453_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_453_inst_req_1;
      ADD_u16_u16_453_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : SLT_i32_u1_409_inst 
    ApIntSlt_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_406_wire & type_cast_408_wire;
      iNsTr_6_410 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_409_inst_req_0;
      SLT_i32_u1_409_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_409_inst_req_1;
      SLT_i32_u1_409_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_1_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : type_cast_424_inst 
    ApIntToApFloatUnsigned_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_9_421;
      iNsTr_10_425 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_424_inst_req_0;
      type_cast_424_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_424_inst_req_1;
      type_cast_424_inst_ack_1 <= ackR_unguarded(0);
      ApIntToApFloatUnsigned_group_2_gI: SplitGuardInterface generic map(name => "ApIntToApFloatUnsigned_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApFloatUnsigned",
          name => "ApIntToApFloatUnsigned_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 8, 
          output_mantissa_width => 23, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : LOAD_ncols_398_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_ncols_398_load_0_req_0;
      LOAD_ncols_398_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ncols_398_load_0_req_1;
      LOAD_ncols_398_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncols_398_word_address_0;
      LOAD_ncols_398_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_447_load_0 ptr_deref_428_load_0 ptr_deref_391_load_0 ptr_deref_420_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_447_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_428_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_391_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_420_load_0_req_0;
      ptr_deref_447_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_428_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_391_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_420_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_447_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_428_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_391_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_420_load_0_req_1;
      ptr_deref_447_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_428_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_391_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_420_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_447_word_address_0 & ptr_deref_428_word_address_0 & ptr_deref_391_word_address_0 & ptr_deref_420_word_address_0;
      ptr_deref_447_data_0 <= data_out(63 downto 48);
      ptr_deref_428_data_0 <= data_out(47 downto 32);
      ptr_deref_391_data_0 <= data_out(31 downto 16);
      ptr_deref_420_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_15_lr_req(0),
          mack => memory_space_15_lr_ack(0),
          maddr => memory_space_15_lr_addr(0 downto 0),
          mtag => memory_space_15_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_15_lc_req(0),
          mack => memory_space_15_lc_ack(0),
          mdata => memory_space_15_lc_data(15 downto 0),
          mtag => memory_space_15_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_456_store_0 ptr_deref_383_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_456_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_383_store_0_req_0;
      ptr_deref_456_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_383_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_456_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_383_store_0_req_1;
      ptr_deref_456_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_383_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_456_word_address_0 & ptr_deref_383_word_address_0;
      data_in <= ptr_deref_456_data_0 & ptr_deref_383_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_15_sr_req(0),
          mack => memory_space_15_sr_ack(0),
          maddr => memory_space_15_sr_addr(0 downto 0),
          mdata => memory_space_15_sr_data(15 downto 0),
          mtag => memory_space_15_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_15_sc_req(0),
          mack => memory_space_15_sc_ack(0),
          mtag => memory_space_15_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_440_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_440_store_0_req_0;
      ptr_deref_440_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_440_store_0_req_1;
      ptr_deref_440_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_440_word_address_0;
      data_in <= ptr_deref_440_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(9 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_15: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_15",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_15_lr_addr,
      lr_req_in => memory_space_15_lr_req,
      lr_ack_out => memory_space_15_lr_ack,
      lr_tag_in => memory_space_15_lr_tag,
      lc_req_in => memory_space_15_lc_req,
      lc_ack_out => memory_space_15_lc_ack,
      lc_data_out => memory_space_15_lc_data,
      lc_tag_out => memory_space_15_lc_tag,
      sr_addr_in => memory_space_15_sr_addr,
      sr_data_in => memory_space_15_sr_data,
      sr_req_in => memory_space_15_sr_req,
      sr_ack_out => memory_space_15_sr_ack,
      sr_tag_in => memory_space_15_sr_tag,
      sc_req_in=> memory_space_15_sc_req,
      sc_ack_out => memory_space_15_sc_ack,
      sc_tag_out => memory_space_15_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end initialize_aPriori_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readCodeBlock is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    code_block_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    code_block_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    code_block_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readCodeBlock;
architecture readCodeBlock_arch of readCodeBlock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal readCodeBlock_CP_2991_start: Boolean;
  signal readCodeBlock_CP_2991_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_479_store_0_req_0 : boolean;
  signal ptr_deref_479_store_0_ack_0 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal SLT_i32_u1_505_inst_req_0 : boolean;
  signal type_cast_491_inst_ack_0 : boolean;
  signal type_cast_491_inst_req_0 : boolean;
  signal type_cast_498_inst_ack_1 : boolean;
  signal type_cast_491_inst_ack_1 : boolean;
  signal SLT_i32_u1_505_inst_ack_0 : boolean;
  signal SLT_i32_u1_505_inst_req_1 : boolean;
  signal SLT_i32_u1_505_inst_ack_1 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal type_cast_498_inst_req_1 : boolean;
  signal type_cast_491_inst_req_1 : boolean;
  signal if_stmt_507_branch_req_0 : boolean;
  signal ptr_deref_487_load_0_ack_1 : boolean;
  signal ptr_deref_487_load_0_req_1 : boolean;
  signal LOAD_ncols_494_load_0_ack_1 : boolean;
  signal ptr_deref_487_load_0_ack_0 : boolean;
  signal ptr_deref_487_load_0_req_0 : boolean;
  signal LOAD_ncols_494_load_0_req_1 : boolean;
  signal LOAD_ncols_494_load_0_ack_0 : boolean;
  signal LOAD_ncols_494_load_0_req_0 : boolean;
  signal ptr_deref_479_store_0_ack_1 : boolean;
  signal ptr_deref_479_store_0_req_1 : boolean;
  signal if_stmt_507_branch_ack_1 : boolean;
  signal if_stmt_507_branch_ack_0 : boolean;
  signal RPIPE_code_block_in_515_inst_req_0 : boolean;
  signal RPIPE_code_block_in_515_inst_ack_0 : boolean;
  signal RPIPE_code_block_in_515_inst_req_1 : boolean;
  signal RPIPE_code_block_in_515_inst_ack_1 : boolean;
  signal ptr_deref_518_store_0_req_0 : boolean;
  signal ptr_deref_518_store_0_ack_0 : boolean;
  signal ptr_deref_518_store_0_req_1 : boolean;
  signal ptr_deref_518_store_0_ack_1 : boolean;
  signal ptr_deref_523_load_0_req_0 : boolean;
  signal ptr_deref_523_load_0_ack_0 : boolean;
  signal ptr_deref_523_load_0_req_1 : boolean;
  signal ptr_deref_523_load_0_ack_1 : boolean;
  signal ptr_deref_527_load_0_req_0 : boolean;
  signal ptr_deref_527_load_0_ack_0 : boolean;
  signal ptr_deref_527_load_0_req_1 : boolean;
  signal ptr_deref_527_load_0_ack_1 : boolean;
  signal type_cast_531_inst_req_0 : boolean;
  signal type_cast_531_inst_ack_0 : boolean;
  signal type_cast_531_inst_req_1 : boolean;
  signal type_cast_531_inst_ack_1 : boolean;
  signal addr_of_536_final_reg_req_0 : boolean;
  signal addr_of_536_final_reg_ack_0 : boolean;
  signal addr_of_536_final_reg_req_1 : boolean;
  signal addr_of_536_final_reg_ack_1 : boolean;
  signal ptr_deref_539_store_0_req_0 : boolean;
  signal ptr_deref_539_store_0_ack_0 : boolean;
  signal ptr_deref_539_store_0_req_1 : boolean;
  signal ptr_deref_539_store_0_ack_1 : boolean;
  signal ptr_deref_546_load_0_req_0 : boolean;
  signal ptr_deref_546_load_0_ack_0 : boolean;
  signal ptr_deref_546_load_0_req_1 : boolean;
  signal ptr_deref_546_load_0_ack_1 : boolean;
  signal ADD_u8_u8_552_inst_req_0 : boolean;
  signal ADD_u8_u8_552_inst_ack_0 : boolean;
  signal ADD_u8_u8_552_inst_req_1 : boolean;
  signal ADD_u8_u8_552_inst_ack_1 : boolean;
  signal ptr_deref_555_store_0_req_0 : boolean;
  signal ptr_deref_555_store_0_ack_0 : boolean;
  signal ptr_deref_555_store_0_req_1 : boolean;
  signal ptr_deref_555_store_0_ack_1 : boolean;
  signal memory_space_16_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_16_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_16_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_16_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_16_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_16_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_17_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_17_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_17_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_17_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_17_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readCodeBlock_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readCodeBlock_CP_2991_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readCodeBlock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readCodeBlock_CP_2991_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readCodeBlock_CP_2991_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readCodeBlock_CP_2991_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readCodeBlock_CP_2991: Block -- control-path 
    signal readCodeBlock_CP_2991_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    readCodeBlock_CP_2991_elements(0) <= readCodeBlock_CP_2991_start;
    readCodeBlock_CP_2991_symbol <= readCodeBlock_CP_2991_elements(81);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_466/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	12 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482__entry__
      -- CP-element group 1: 	 branch_block_stmt_466/branch_block_stmt_466__entry__
      -- 
    readCodeBlock_CP_2991_elements(1) <= readCodeBlock_CP_2991_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	14 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	65 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_466/bb_0_bb_1
      -- CP-element group 2: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482__exit__
      -- 
    readCodeBlock_CP_2991_elements(2) <= readCodeBlock_CP_2991_elements(14);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	68 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	15 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506__entry__
      -- CP-element group 3: 	 branch_block_stmt_466/merge_stmt_484__exit__
      -- 
    readCodeBlock_CP_2991_elements(3) <= readCodeBlock_CP_2991_elements(68);
    -- CP-element group 4:  branch  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	26 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4: 	28 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_466/if_stmt_507__entry__
      -- CP-element group 4: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506__exit__
      -- 
    readCodeBlock_CP_2991_elements(4) <= readCodeBlock_CP_2991_elements(26);
    -- CP-element group 5:  merge  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	36 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_466/assign_stmt_516__entry__
      -- CP-element group 5: 	 branch_block_stmt_466/merge_stmt_513__exit__
      -- 
    readCodeBlock_CP_2991_elements(5) <= readCodeBlock_CP_2991_elements(71);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	38 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	39 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541__entry__
      -- CP-element group 6: 	 branch_block_stmt_466/assign_stmt_516__exit__
      -- 
    readCodeBlock_CP_2991_elements(6) <= readCodeBlock_CP_2991_elements(38);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	55 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	72 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_466/bb_2_bb_3
      -- CP-element group 7: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541__exit__
      -- 
    readCodeBlock_CP_2991_elements(7) <= readCodeBlock_CP_2991_elements(55);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	74 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	56 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557__entry__
      -- CP-element group 8: 	 branch_block_stmt_466/merge_stmt_543__exit__
      -- 
    readCodeBlock_CP_2991_elements(8) <= readCodeBlock_CP_2991_elements(74);
    -- CP-element group 9:  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	63 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	66 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_466/bb_3_bb_1
      -- CP-element group 9: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557__exit__
      -- 
    readCodeBlock_CP_2991_elements(9) <= readCodeBlock_CP_2991_elements(63);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	77 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	78 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_466/return__
      -- CP-element group 10: 	 branch_block_stmt_466/merge_stmt_559__exit__
      -- 
    readCodeBlock_CP_2991_elements(10) <= readCodeBlock_CP_2991_elements(77);
    -- CP-element group 11:  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	80 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	81 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_466/merge_stmt_561__exit__
      -- CP-element group 11: 	 branch_block_stmt_466/branch_block_stmt_466__exit__
      -- 
    readCodeBlock_CP_2991_elements(11) <= readCodeBlock_CP_2991_elements(80);
    -- CP-element group 12:  fork  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	1 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (31) 
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_word_address_calculated
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_addr_resize/$exit
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_word_addrgen/root_register_ack
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/ptr_deref_479_Split/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_word_addrgen/$exit
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/word_0/rr
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_address_resized
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_addr_resize/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_update_start_
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_word_addrgen/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/word_0/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_plus_offset/sum_rename_ack
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_root_address_calculated
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/ptr_deref_479_Split/$exit
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/word_0/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_address_calculated
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_addr_resize/base_resize_ack
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/ptr_deref_479_Split/split_ack
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_plus_offset/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_plus_offset/$exit
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_base_addr_resize/base_resize_req
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/$entry
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_word_addrgen/root_register_req
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/word_0/cr
      -- CP-element group 12: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/ptr_deref_479_Split/split_req
      -- 
    cr_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(12), ack => ptr_deref_479_store_0_req_1); -- 
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(12), ack => ptr_deref_479_store_0_req_0); -- 
    readCodeBlock_CP_2991_elements(12) <= readCodeBlock_CP_2991_elements(1);
    -- CP-element group 13:  transition  input  no-bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_sample_completed_
      -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_store_0_ack_0, ack => readCodeBlock_CP_2991_elements(13)); -- 
    -- CP-element group 14:  transition  input  no-bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	2 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/$exit
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_466/assign_stmt_473_to_assign_stmt_482/ptr_deref_479_Update/word_access_complete/word_0/$exit
      -- 
    ca_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_store_0_ack_1, ack => readCodeBlock_CP_2991_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	26 
    -- CP-element group 15:  members (48) 
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_update_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_update_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_update_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_update_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/word_0/cr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/word_0/cr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_addr_resize/base_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_addr_resize/base_resize_req
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_addr_resize/$exit
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_addr_resize/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_address_resized
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_base_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_update_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/$entry
      -- 
    cr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => ptr_deref_487_load_0_req_1); -- 
    rr_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => ptr_deref_487_load_0_req_0); -- 
    cr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => type_cast_491_inst_req_1); -- 
    cr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => LOAD_ncols_494_load_0_req_1); -- 
    rr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => LOAD_ncols_494_load_0_req_0); -- 
    cr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => type_cast_498_inst_req_1); -- 
    cr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(15), ack => SLT_i32_u1_505_inst_req_1); -- 
    readCodeBlock_CP_2991_elements(15) <= readCodeBlock_CP_2991_elements(3);
    -- CP-element group 16:  transition  input  no-bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/word_0/ra
      -- CP-element group 16: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_sample_completed_
      -- 
    ra_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_487_load_0_ack_0, ack => readCodeBlock_CP_2991_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  no-bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (12) 
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/ptr_deref_487_Merge/merge_ack
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/ptr_deref_487_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/ptr_deref_487_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/ptr_deref_487_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/ptr_deref_487_update_completed_
      -- 
    ca_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_487_load_0_ack_1, ack => readCodeBlock_CP_2991_elements(17)); -- 
    rr_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(17), ack => type_cast_491_inst_req_0); -- 
    -- CP-element group 18:  transition  input  no-bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_sample_completed_
      -- 
    ra_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_0, ack => readCodeBlock_CP_2991_elements(18)); -- 
    -- CP-element group 19:  transition  input  no-bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_491_update_completed_
      -- 
    ca_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_491_inst_ack_1, ack => readCodeBlock_CP_2991_elements(19)); -- 
    -- CP-element group 20:  transition  input  no-bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/word_0/ra
      -- CP-element group 20: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Sample/$exit
      -- 
    ra_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_494_load_0_ack_0, ack => readCodeBlock_CP_2991_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  no-bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (12) 
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/LOAD_ncols_494_Merge/merge_ack
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/LOAD_ncols_494_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/LOAD_ncols_494_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/LOAD_ncols_494_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/LOAD_ncols_494_Update/$exit
      -- 
    ca_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_494_load_0_ack_1, ack => readCodeBlock_CP_2991_elements(21)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(21), ack => type_cast_498_inst_req_0); -- 
    -- CP-element group 22:  transition  input  no-bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Sample/$exit
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_0, ack => readCodeBlock_CP_2991_elements(22)); -- 
    -- CP-element group 23:  transition  input  no-bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/type_cast_498_Update/ca
      -- 
    ca_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_1, ack => readCodeBlock_CP_2991_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_sample_start_
      -- 
    rr_3195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(24), ack => SLT_i32_u1_505_inst_req_0); -- 
    readCodeBlock_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "readCodeBlock_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readCodeBlock_CP_2991_elements(19) & readCodeBlock_CP_2991_elements(23);
      gj_readCodeBlock_cp_element_group_24 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readCodeBlock_CP_2991_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  no-bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_sample_completed_
      -- 
    ra_3196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_505_inst_ack_0, ack => readCodeBlock_CP_2991_elements(25)); -- 
    -- CP-element group 26:  transition  input  no-bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	4 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/SLT_i32_u1_505_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_466/assign_stmt_488_to_assign_stmt_506/$exit
      -- 
    ca_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_505_inst_ack_1, ack => readCodeBlock_CP_2991_elements(26)); -- 
    -- CP-element group 27:  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_466/if_stmt_507_dead_link/$entry
      -- 
    readCodeBlock_CP_2991_elements(27) <= readCodeBlock_CP_2991_elements(4);
    -- CP-element group 28:  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	4 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_466/if_stmt_507_eval_test/$entry
      -- CP-element group 28: 	 branch_block_stmt_466/if_stmt_507_eval_test/$exit
      -- CP-element group 28: 	 branch_block_stmt_466/if_stmt_507_eval_test/branch_req
      -- 
    branch_req_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(28), ack => if_stmt_507_branch_req_0); -- 
    readCodeBlock_CP_2991_elements(28) <= readCodeBlock_CP_2991_elements(4);
    -- CP-element group 29:  branch  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_466/R_iNsTr_6_508_place
      -- 
    readCodeBlock_CP_2991_elements(29) <= readCodeBlock_CP_2991_elements(28);
    -- CP-element group 30:  transition  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_466/if_stmt_507_if_link/$entry
      -- 
    readCodeBlock_CP_2991_elements(30) <= readCodeBlock_CP_2991_elements(29);
    -- CP-element group 31:  transition  input  no-bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_466/if_stmt_507_if_link/$exit
      -- CP-element group 31: 	 branch_block_stmt_466/if_stmt_507_if_link/if_choice_transition
      -- 
    if_choice_transition_3214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_507_branch_ack_1, ack => readCodeBlock_CP_2991_elements(31)); -- 
    -- CP-element group 32:  transition  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_466/if_stmt_507_else_link/$entry
      -- 
    readCodeBlock_CP_2991_elements(32) <= readCodeBlock_CP_2991_elements(29);
    -- CP-element group 33:  transition  input  no-bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_466/if_stmt_507_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_466/if_stmt_507_else_link/else_choice_transition
      -- 
    else_choice_transition_3218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_507_branch_ack_0, ack => readCodeBlock_CP_2991_elements(33)); -- 
    -- CP-element group 34:  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	69 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_466/bb_1_bb_2
      -- 
    readCodeBlock_CP_2991_elements(34) <= readCodeBlock_CP_2991_elements(31);
    -- CP-element group 35:  place  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	75 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_466/bb_1_bb_4
      -- 
    readCodeBlock_CP_2991_elements(35) <= readCodeBlock_CP_2991_elements(33);
    -- CP-element group 36:  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	5 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_466/assign_stmt_516/$entry
      -- CP-element group 36: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Sample/rr
      -- 
    rr_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(36), ack => RPIPE_code_block_in_515_inst_req_0); -- 
    readCodeBlock_CP_2991_elements(36) <= readCodeBlock_CP_2991_elements(5);
    -- CP-element group 37:  transition  input  output  no-bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_update_start_
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Update/cr
      -- 
    ra_3232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_code_block_in_515_inst_ack_0, ack => readCodeBlock_CP_2991_elements(37)); -- 
    cr_3236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(37), ack => RPIPE_code_block_in_515_inst_req_1); -- 
    -- CP-element group 38:  transition  input  no-bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	6 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_466/assign_stmt_516/$exit
      -- CP-element group 38: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_466/assign_stmt_516/RPIPE_code_block_in_515_Update/ca
      -- 
    ca_3237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_code_block_in_515_inst_ack_1, ack => readCodeBlock_CP_2991_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	6 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	42 
    -- CP-element group 39: 	44 
    -- CP-element group 39: 	45 
    -- CP-element group 39: 	46 
    -- CP-element group 39: 	48 
    -- CP-element group 39: 	50 
    -- CP-element group 39: 	53 
    -- CP-element group 39:  members (89) 
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/ptr_deref_518_Split/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/ptr_deref_518_Split/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/ptr_deref_518_Split/split_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/ptr_deref_518_Split/split_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/word_0/rr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/word_0/rr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_complete/req
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_update_start_
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/word_0/cr
      -- 
    cr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_518_store_0_req_1); -- 
    rr_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_518_store_0_req_0); -- 
    cr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_523_load_0_req_1); -- 
    cr_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_527_load_0_req_1); -- 
    rr_3373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_527_load_0_req_0); -- 
    cr_3403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => type_cast_531_inst_req_1); -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => addr_of_536_final_reg_req_1); -- 
    cr_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(39), ack => ptr_deref_539_store_0_req_1); -- 
    readCodeBlock_CP_2991_elements(39) <= readCodeBlock_CP_2991_elements(6);
    -- CP-element group 40:  transition  input  no-bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	54 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Sample/word_access_start/word_0/ra
      -- 
    ra_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_518_store_0_ack_0, ack => readCodeBlock_CP_2991_elements(40)); -- 
    -- CP-element group 41:  transition  input  no-bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	55 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_Update/word_access_complete/word_0/ca
      -- 
    ca_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_518_store_0_ack_1, ack => readCodeBlock_CP_2991_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: 	54 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/word_0/rr
      -- 
    rr_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(42), ack => ptr_deref_523_load_0_req_0); -- 
    readCodeBlock_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "readCodeBlock_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readCodeBlock_CP_2991_elements(39) & readCodeBlock_CP_2991_elements(54);
      gj_readCodeBlock_cp_element_group_42 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readCodeBlock_CP_2991_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  no-bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Sample/word_access_start/word_0/ra
      -- 
    ra_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_523_load_0_ack_0, ack => readCodeBlock_CP_2991_elements(43)); -- 
    -- CP-element group 44:  transition  input  no-bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	39 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/ptr_deref_523_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/ptr_deref_523_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/ptr_deref_523_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_523_Update/ptr_deref_523_Merge/merge_ack
      -- 
    ca_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_523_load_0_ack_1, ack => readCodeBlock_CP_2991_elements(44)); -- 
    -- CP-element group 45:  transition  input  no-bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	39 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Sample/word_access_start/word_0/ra
      -- 
    ra_3374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_527_load_0_ack_0, ack => readCodeBlock_CP_2991_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  no-bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	39 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (12) 
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/ptr_deref_527_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/ptr_deref_527_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/ptr_deref_527_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_527_Update/ptr_deref_527_Merge/merge_ack
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Sample/rr
      -- 
    ca_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_527_load_0_ack_1, ack => readCodeBlock_CP_2991_elements(46)); -- 
    rr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(46), ack => type_cast_531_inst_req_0); -- 
    -- CP-element group 47:  transition  input  no-bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Sample/ra
      -- 
    ra_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_0, ack => readCodeBlock_CP_2991_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  no-bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	39 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (27) 
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/type_cast_531_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_resized_0
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_scaled_0
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_computed_0
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_resize_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_resize_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_resize_0/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_resize_0/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_scale_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_scale_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_scale_0/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_index_scale_0/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_final_index_sum_regn/$entry
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_final_index_sum_regn/$exit
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_final_index_sum_regn/req
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_final_index_sum_regn/ack
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/array_obj_ref_535_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_request/req
      -- 
    ca_3404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_1, ack => readCodeBlock_CP_2991_elements(48)); -- 
    req_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(48), ack => addr_of_536_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  no-bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	55 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_request/ack
      -- 
    ack_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_536_final_reg_ack_0, ack => readCodeBlock_CP_2991_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  no-bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	39 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/addr_of_536_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_word_addrgen/root_register_ack
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_536_final_reg_ack_1, ack => readCodeBlock_CP_2991_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/ptr_deref_539_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/ptr_deref_539_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/ptr_deref_539_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/ptr_deref_539_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/word_0/rr
      -- 
    rr_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(51), ack => ptr_deref_539_store_0_req_0); -- 
    readCodeBlock_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "readCodeBlock_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readCodeBlock_CP_2991_elements(44) & readCodeBlock_CP_2991_elements(50);
      gj_readCodeBlock_cp_element_group_51 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readCodeBlock_CP_2991_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  no-bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Sample/word_access_start/word_0/ra
      -- 
    ra_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_539_store_0_ack_0, ack => readCodeBlock_CP_2991_elements(52)); -- 
    -- CP-element group 53:  transition  input  no-bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	39 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_539_Update/word_access_complete/word_0/ca
      -- 
    ca_3493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_539_store_0_ack_1, ack => readCodeBlock_CP_2991_elements(53)); -- 
    -- CP-element group 54:  transition  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	40 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	42 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/ptr_deref_518_ptr_deref_523_delay
      -- 
    -- Element group readCodeBlock_CP_2991_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => readCodeBlock_CP_2991_elements(40), ack => readCodeBlock_CP_2991_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  join  transition  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	41 
    -- CP-element group 55: 	49 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	7 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_466/assign_stmt_520_to_assign_stmt_541/$exit
      -- 
    readCodeBlock_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "readCodeBlock_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readCodeBlock_CP_2991_elements(41) & readCodeBlock_CP_2991_elements(49) & readCodeBlock_CP_2991_elements(53);
      gj_readCodeBlock_cp_element_group_55 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readCodeBlock_CP_2991_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	8 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	61 
    -- CP-element group 56: 	63 
    -- CP-element group 56:  members (51) 
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_update_start_
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_update_start_
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_update_start_
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/word_0/cr
      -- 
    cr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(56), ack => ptr_deref_546_load_0_req_1); -- 
    rr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(56), ack => ptr_deref_546_load_0_req_0); -- 
    cr_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(56), ack => ADD_u8_u8_552_inst_req_1); -- 
    cr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(56), ack => ptr_deref_555_store_0_req_1); -- 
    readCodeBlock_CP_2991_elements(56) <= readCodeBlock_CP_2991_elements(8);
    -- CP-element group 57:  transition  input  no-bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	64 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/$exit
      -- CP-element group 57: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Sample/word_access_start/word_0/ra
      -- 
    ra_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_546_load_0_ack_0, ack => readCodeBlock_CP_2991_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  no-bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (12) 
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/word_access_complete/word_0/ca
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/ptr_deref_546_Merge/$entry
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/ptr_deref_546_Merge/$exit
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/ptr_deref_546_Merge/merge_req
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_Update/ptr_deref_546_Merge/merge_ack
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Sample/rr
      -- 
    ca_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_546_load_0_ack_1, ack => readCodeBlock_CP_2991_elements(58)); -- 
    rr_3555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(58), ack => ADD_u8_u8_552_inst_req_0); -- 
    -- CP-element group 59:  transition  input  no-bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Sample/ra
      -- 
    ra_3556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_552_inst_ack_0, ack => readCodeBlock_CP_2991_elements(59)); -- 
    -- CP-element group 60:  transition  input  no-bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ADD_u8_u8_552_Update/ca
      -- 
    ca_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_552_inst_ack_1, ack => readCodeBlock_CP_2991_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  no-bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	56 
    -- CP-element group 61: 	60 
    -- CP-element group 61: 	64 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/ptr_deref_555_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/ptr_deref_555_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/ptr_deref_555_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/ptr_deref_555_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/word_0/rr
      -- 
    rr_3599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readCodeBlock_CP_2991_elements(61), ack => ptr_deref_555_store_0_req_0); -- 
    readCodeBlock_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 33) := "readCodeBlock_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readCodeBlock_CP_2991_elements(56) & readCodeBlock_CP_2991_elements(60) & readCodeBlock_CP_2991_elements(64);
      gj_readCodeBlock_cp_element_group_61 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readCodeBlock_CP_2991_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  no-bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Sample/word_access_start/word_0/ra
      -- 
    ra_3600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_555_store_0_ack_0, ack => readCodeBlock_CP_2991_elements(62)); -- 
    -- CP-element group 63:  transition  input  no-bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	56 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	9 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/$exit
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_555_Update/word_access_complete/word_0/ca
      -- 
    ca_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_555_store_0_ack_1, ack => readCodeBlock_CP_2991_elements(63)); -- 
    -- CP-element group 64:  transition  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	57 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	61 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_466/assign_stmt_547_to_assign_stmt_557/ptr_deref_546_ptr_deref_555_delay
      -- 
    -- Element group readCodeBlock_CP_2991_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => readCodeBlock_CP_2991_elements(57), ack => readCodeBlock_CP_2991_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  transition  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	2 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_466/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_466/bb_0_bb_1_PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(65) <= readCodeBlock_CP_2991_elements(2);
    -- CP-element group 66:  transition  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	9 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_466/bb_3_bb_1_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_466/bb_3_bb_1_PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(66) <= readCodeBlock_CP_2991_elements(9);
    -- CP-element group 67:  merge  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_466/merge_stmt_484_PhiReqMerge
      -- 
    readCodeBlock_CP_2991_elements(67) <= OrReduce(readCodeBlock_CP_2991_elements(65) & readCodeBlock_CP_2991_elements(66));
    -- CP-element group 68:  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	3 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_466/merge_stmt_484_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_466/merge_stmt_484_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_466/merge_stmt_484_PhiAck/dummy
      -- 
    readCodeBlock_CP_2991_elements(68) <= readCodeBlock_CP_2991_elements(67);
    -- CP-element group 69:  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	34 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_466/bb_1_bb_2_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_466/bb_1_bb_2_PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(69) <= readCodeBlock_CP_2991_elements(34);
    -- CP-element group 70:  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_466/merge_stmt_513_PhiReqMerge
      -- 
    readCodeBlock_CP_2991_elements(70) <= readCodeBlock_CP_2991_elements(69);
    -- CP-element group 71:  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	5 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_466/merge_stmt_513_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_466/merge_stmt_513_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_466/merge_stmt_513_PhiAck/dummy
      -- 
    readCodeBlock_CP_2991_elements(71) <= readCodeBlock_CP_2991_elements(70);
    -- CP-element group 72:  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	7 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_466/bb_2_bb_3_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_466/bb_2_bb_3_PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(72) <= readCodeBlock_CP_2991_elements(7);
    -- CP-element group 73:  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_466/merge_stmt_543_PhiReqMerge
      -- 
    readCodeBlock_CP_2991_elements(73) <= readCodeBlock_CP_2991_elements(72);
    -- CP-element group 74:  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	8 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_466/merge_stmt_543_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_466/merge_stmt_543_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_466/merge_stmt_543_PhiAck/dummy
      -- 
    readCodeBlock_CP_2991_elements(74) <= readCodeBlock_CP_2991_elements(73);
    -- CP-element group 75:  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	35 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_466/bb_1_bb_4_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_466/bb_1_bb_4_PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(75) <= readCodeBlock_CP_2991_elements(35);
    -- CP-element group 76:  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_466/merge_stmt_559_PhiReqMerge
      -- 
    readCodeBlock_CP_2991_elements(76) <= readCodeBlock_CP_2991_elements(75);
    -- CP-element group 77:  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	10 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_466/merge_stmt_559_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_466/merge_stmt_559_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_466/merge_stmt_559_PhiAck/dummy
      -- 
    readCodeBlock_CP_2991_elements(77) <= readCodeBlock_CP_2991_elements(76);
    -- CP-element group 78:  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	10 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_466/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_466/return___PhiReq/$exit
      -- 
    readCodeBlock_CP_2991_elements(78) <= readCodeBlock_CP_2991_elements(10);
    -- CP-element group 79:  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_466/merge_stmt_561_PhiReqMerge
      -- 
    readCodeBlock_CP_2991_elements(79) <= readCodeBlock_CP_2991_elements(78);
    -- CP-element group 80:  transition  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	11 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_466/merge_stmt_561_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_466/merge_stmt_561_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_466/merge_stmt_561_PhiAck/dummy
      -- 
    readCodeBlock_CP_2991_elements(80) <= readCodeBlock_CP_2991_elements(79);
    -- CP-element group 81:  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	11 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_466/$exit
      -- CP-element group 81: 	 $exit
      -- 
    readCodeBlock_CP_2991_elements(81) <= readCodeBlock_CP_2991_elements(11);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_473 : std_logic_vector(31 downto 0);
    signal LOAD_ncols_494_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_494_word_address_0 : std_logic_vector(0 downto 0);
    signal R_iNsTr_14_534_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_14_534_scaled : std_logic_vector(9 downto 0);
    signal array_obj_ref_535_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_535_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_535_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_535_root_address : std_logic_vector(9 downto 0);
    signal code_bit_477 : std_logic_vector(31 downto 0);
    signal iNsTr_10_516 : std_logic_vector(31 downto 0);
    signal iNsTr_12_524 : std_logic_vector(31 downto 0);
    signal iNsTr_13_528 : std_logic_vector(7 downto 0);
    signal iNsTr_14_532 : std_logic_vector(63 downto 0);
    signal iNsTr_15_537 : std_logic_vector(31 downto 0);
    signal iNsTr_19_547 : std_logic_vector(7 downto 0);
    signal iNsTr_20_553 : std_logic_vector(7 downto 0);
    signal iNsTr_2_488 : std_logic_vector(7 downto 0);
    signal iNsTr_3_492 : std_logic_vector(31 downto 0);
    signal iNsTr_4_495 : std_logic_vector(15 downto 0);
    signal iNsTr_5_499 : std_logic_vector(31 downto 0);
    signal iNsTr_6_506 : std_logic_vector(0 downto 0);
    signal ptr_deref_479_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_479_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_479_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_479_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_479_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_479_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_487_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_487_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_487_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_487_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_487_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_518_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_518_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_518_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_518_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_518_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_518_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_523_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_523_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_523_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_523_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_523_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_527_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_527_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_527_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_527_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_527_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_539_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_539_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_539_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_539_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_539_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_539_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_546_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_546_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_546_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_546_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_546_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_555_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_555_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_555_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_555_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_555_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_555_word_offset_0 : std_logic_vector(0 downto 0);
    signal type_cast_481_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_502_wire : std_logic_vector(31 downto 0);
    signal type_cast_504_wire : std_logic_vector(31 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(7 downto 0);
    signal xxreadCodeBlockxxbodyxxI_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxreadCodeBlockxxbodyxxcode_bit_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    I_473 <= "00000000000000000000000000000000";
    LOAD_ncols_494_word_address_0 <= "0";
    array_obj_ref_535_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_535_resized_base_address <= "0000000000";
    code_bit_477 <= "00000000000000000000000000000000";
    ptr_deref_479_word_offset_0 <= "0";
    ptr_deref_487_word_offset_0 <= "0";
    ptr_deref_518_word_offset_0 <= "0";
    ptr_deref_523_word_offset_0 <= "0";
    ptr_deref_527_word_offset_0 <= "0";
    ptr_deref_539_word_offset_0 <= "0000000000";
    ptr_deref_546_word_offset_0 <= "0";
    ptr_deref_555_word_offset_0 <= "0";
    type_cast_481_wire_constant <= "00000000";
    type_cast_551_wire_constant <= "00000001";
    xxreadCodeBlockxxbodyxxI_alloc_base_address <= "0";
    xxreadCodeBlockxxbodyxxcode_bit_alloc_base_address <= "0";
    addr_of_536_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_536_final_reg_req_0;
      addr_of_536_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_536_final_reg_req_1;
      addr_of_536_final_reg_ack_1<= rack(0);
      addr_of_536_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_536_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_535_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_15_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_491_inst_req_0;
      type_cast_491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_491_inst_req_1;
      type_cast_491_inst_ack_1<= rack(0);
      type_cast_491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_2_488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_3_492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_498_inst_req_0;
      type_cast_498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_498_inst_req_1;
      type_cast_498_inst_ack_1<= rack(0);
      type_cast_498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_4_495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_5_499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_502_inst
    process(iNsTr_3_492) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_3_492(31 downto 0);
      type_cast_502_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_504_inst
    process(iNsTr_5_499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_5_499(31 downto 0);
      type_cast_504_wire <= tmp_var; -- 
    end process;
    type_cast_531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_531_inst_req_0;
      type_cast_531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_531_inst_req_1;
      type_cast_531_inst_ack_1<= rack(0);
      type_cast_531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_13_528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_ncols_494_gather_scatter
    process(LOAD_ncols_494_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_494_data_0;
      ov(15 downto 0) := iv;
      iNsTr_4_495 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_535_index_0_rename
    process(R_iNsTr_14_534_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_14_534_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_14_534_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_535_index_0_resize
    process(iNsTr_14_532) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_14_532;
      ov := iv(9 downto 0);
      R_iNsTr_14_534_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_535_index_offset
    process(R_iNsTr_14_534_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_14_534_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_535_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_535_root_address_inst
    process(array_obj_ref_535_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_535_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_535_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_addr_0
    process(ptr_deref_479_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_479_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_base_resize
    process(I_473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_473;
      ov := iv(0 downto 0);
      ptr_deref_479_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_gather_scatter
    process(type_cast_481_wire_constant) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_481_wire_constant;
      ov(7 downto 0) := iv;
      ptr_deref_479_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_root_address_inst
    process(ptr_deref_479_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_479_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_addr_0
    process(ptr_deref_487_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_487_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_487_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_base_resize
    process(I_473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_473;
      ov := iv(0 downto 0);
      ptr_deref_487_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_gather_scatter
    process(ptr_deref_487_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_487_data_0;
      ov(7 downto 0) := iv;
      iNsTr_2_488 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_root_address_inst
    process(ptr_deref_487_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_487_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_487_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_addr_0
    process(ptr_deref_518_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_518_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_518_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_base_resize
    process(code_bit_477) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := code_bit_477;
      ov := iv(0 downto 0);
      ptr_deref_518_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_gather_scatter
    process(iNsTr_10_516) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_516;
      ov(31 downto 0) := iv;
      ptr_deref_518_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_518_root_address_inst
    process(ptr_deref_518_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_518_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_518_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_addr_0
    process(ptr_deref_523_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_523_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_523_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_base_resize
    process(code_bit_477) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := code_bit_477;
      ov := iv(0 downto 0);
      ptr_deref_523_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_gather_scatter
    process(ptr_deref_523_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_523_data_0;
      ov(31 downto 0) := iv;
      iNsTr_12_524 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_523_root_address_inst
    process(ptr_deref_523_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_523_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_523_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_527_addr_0
    process(ptr_deref_527_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_527_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_527_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_527_base_resize
    process(I_473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_473;
      ov := iv(0 downto 0);
      ptr_deref_527_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_527_gather_scatter
    process(ptr_deref_527_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_527_data_0;
      ov(7 downto 0) := iv;
      iNsTr_13_528 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_527_root_address_inst
    process(ptr_deref_527_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_527_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_527_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_539_addr_0
    process(ptr_deref_539_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_539_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_539_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_539_base_resize
    process(iNsTr_15_537) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_537;
      ov := iv(9 downto 0);
      ptr_deref_539_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_539_gather_scatter
    process(iNsTr_12_524) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_12_524;
      ov(31 downto 0) := iv;
      ptr_deref_539_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_539_root_address_inst
    process(ptr_deref_539_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_539_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_539_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_546_addr_0
    process(ptr_deref_546_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_546_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_546_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_546_base_resize
    process(I_473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_473;
      ov := iv(0 downto 0);
      ptr_deref_546_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_546_gather_scatter
    process(ptr_deref_546_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_546_data_0;
      ov(7 downto 0) := iv;
      iNsTr_19_547 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_546_root_address_inst
    process(ptr_deref_546_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_546_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_546_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_555_addr_0
    process(ptr_deref_555_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_555_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_555_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_555_base_resize
    process(I_473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_473;
      ov := iv(0 downto 0);
      ptr_deref_555_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_555_gather_scatter
    process(iNsTr_20_553) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_20_553;
      ov(7 downto 0) := iv;
      ptr_deref_555_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_555_root_address_inst
    process(ptr_deref_555_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_555_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_555_root_address <= ov(0 downto 0);
      --
    end process;
    if_stmt_507_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_6_506;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_507_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_507_branch_req_0,
          ack0 => if_stmt_507_branch_ack_0,
          ack1 => if_stmt_507_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u8_u8_552_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_19_547;
      iNsTr_20_553 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_552_inst_req_0;
      ADD_u8_u8_552_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_552_inst_req_1;
      ADD_u8_u8_552_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : SLT_i32_u1_505_inst 
    ApIntSlt_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_502_wire & type_cast_504_wire;
      iNsTr_6_506 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_505_inst_req_0;
      SLT_i32_u1_505_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_505_inst_req_1;
      SLT_i32_u1_505_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_1_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared load operator group (0) : LOAD_ncols_494_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_ncols_494_load_0_req_0;
      LOAD_ncols_494_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ncols_494_load_0_req_1;
      LOAD_ncols_494_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncols_494_word_address_0;
      LOAD_ncols_494_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_527_load_0 ptr_deref_487_load_0 ptr_deref_546_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_527_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_487_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_546_load_0_req_0;
      ptr_deref_527_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_487_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_546_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_527_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_487_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_546_load_0_req_1;
      ptr_deref_527_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_487_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_546_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_527_word_address_0 & ptr_deref_487_word_address_0 & ptr_deref_546_word_address_0;
      ptr_deref_527_data_0 <= data_out(23 downto 16);
      ptr_deref_487_data_0 <= data_out(15 downto 8);
      ptr_deref_546_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_16_lr_req(0),
          mack => memory_space_16_lr_ack(0),
          maddr => memory_space_16_lr_addr(0 downto 0),
          mtag => memory_space_16_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_16_lc_req(0),
          mack => memory_space_16_lc_ack(0),
          mdata => memory_space_16_lc_data(7 downto 0),
          mtag => memory_space_16_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_523_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_523_load_0_req_0;
      ptr_deref_523_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_523_load_0_req_1;
      ptr_deref_523_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_523_word_address_0;
      ptr_deref_523_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_17_lr_req(0),
          mack => memory_space_17_lr_ack(0),
          maddr => memory_space_17_lr_addr(0 downto 0),
          mtag => memory_space_17_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_17_lc_req(0),
          mack => memory_space_17_lc_ack(0),
          mdata => memory_space_17_lc_data(31 downto 0),
          mtag => memory_space_17_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_479_store_0 ptr_deref_555_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_479_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_555_store_0_req_0;
      ptr_deref_479_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_555_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_479_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_555_store_0_req_1;
      ptr_deref_479_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_555_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_479_word_address_0 & ptr_deref_555_word_address_0;
      data_in <= ptr_deref_479_data_0 & ptr_deref_555_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_16_sr_req(0),
          mack => memory_space_16_sr_ack(0),
          maddr => memory_space_16_sr_addr(0 downto 0),
          mdata => memory_space_16_sr_data(7 downto 0),
          mtag => memory_space_16_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_16_sc_req(0),
          mack => memory_space_16_sc_ack(0),
          mtag => memory_space_16_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_518_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_518_store_0_req_0;
      ptr_deref_518_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_518_store_0_req_1;
      ptr_deref_518_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_518_word_address_0;
      data_in <= ptr_deref_518_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_17_sr_req(0),
          mack => memory_space_17_sr_ack(0),
          maddr => memory_space_17_sr_addr(0 downto 0),
          mdata => memory_space_17_sr_data(31 downto 0),
          mtag => memory_space_17_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_17_sc_req(0),
          mack => memory_space_17_sc_ack(0),
          mtag => memory_space_17_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_539_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_539_store_0_req_0;
      ptr_deref_539_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_539_store_0_req_1;
      ptr_deref_539_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_539_word_address_0;
      data_in <= ptr_deref_539_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(9 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_code_block_in_515_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_code_block_in_515_inst_req_0;
      RPIPE_code_block_in_515_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_code_block_in_515_inst_req_1;
      RPIPE_code_block_in_515_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_10_516 <= data_out(31 downto 0);
      code_block_in_read_0_gI: SplitGuardInterface generic map(name => "code_block_in_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      code_block_in_read_0: InputPortRevised -- 
        generic map ( name => "code_block_in_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => code_block_in_pipe_read_req(0),
          oack => code_block_in_pipe_read_ack(0),
          odata => code_block_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_16: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_16",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_16_lr_addr,
      lr_req_in => memory_space_16_lr_req,
      lr_ack_out => memory_space_16_lr_ack,
      lr_tag_in => memory_space_16_lr_tag,
      lc_req_in => memory_space_16_lc_req,
      lc_ack_out => memory_space_16_lc_ack,
      lc_data_out => memory_space_16_lc_data,
      lc_tag_out => memory_space_16_lc_tag,
      sr_addr_in => memory_space_16_sr_addr,
      sr_data_in => memory_space_16_sr_data,
      sr_req_in => memory_space_16_sr_req,
      sr_ack_out => memory_space_16_sr_ack,
      sr_tag_in => memory_space_16_sr_tag,
      sc_req_in=> memory_space_16_sc_req,
      sc_ack_out => memory_space_16_sc_ack,
      sc_tag_out => memory_space_16_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_17: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_17",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_17_lr_addr,
      lr_req_in => memory_space_17_lr_req,
      lr_ack_out => memory_space_17_lr_ack,
      lr_tag_in => memory_space_17_lr_tag,
      lc_req_in => memory_space_17_lc_req,
      lc_ack_out => memory_space_17_lc_ack,
      lc_data_out => memory_space_17_lc_data,
      lc_tag_out => memory_space_17_lc_tag,
      sr_addr_in => memory_space_17_sr_addr,
      sr_data_in => memory_space_17_sr_data,
      sr_req_in => memory_space_17_sr_req,
      sr_ack_out => memory_space_17_sr_ack,
      sr_tag_in => memory_space_17_sr_tag,
      sc_req_in=> memory_space_17_sc_req,
      sc_ack_out => memory_space_17_sc_ack,
      sc_tag_out => memory_space_17_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end readCodeBlock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity send_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(31 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    aPriori_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    aPriori_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    aPriori_out_pipe_write_data : out  std_logic_vector(31 downto 0);
    code_block_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    code_block_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    code_block_out_pipe_write_data : out  std_logic_vector(31 downto 0);
    mem_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    mem_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    mem_out_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity send_output;
architecture send_output_arch of send_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(31 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal send_output_CP_3660_start: Boolean;
  signal send_output_CP_3660_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_593_store_0_ack_1 : boolean;
  signal ptr_deref_593_store_0_req_1 : boolean;
  signal ptr_deref_666_load_0_req_0 : boolean;
  signal ptr_deref_593_store_0_req_0 : boolean;
  signal ptr_deref_593_store_0_ack_0 : boolean;
  signal ptr_deref_661_store_0_ack_1 : boolean;
  signal ptr_deref_666_load_0_ack_0 : boolean;
  signal ptr_deref_661_store_0_req_1 : boolean;
  signal ptr_deref_601_load_0_req_0 : boolean;
  signal ptr_deref_601_load_0_ack_0 : boolean;
  signal ptr_deref_601_load_0_req_1 : boolean;
  signal ptr_deref_601_load_0_ack_1 : boolean;
  signal LOAD_nrows_604_load_0_req_0 : boolean;
  signal LOAD_nrows_604_load_0_ack_0 : boolean;
  signal LOAD_nrows_604_load_0_req_1 : boolean;
  signal LOAD_nrows_604_load_0_ack_1 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal ptr_deref_816_load_0_req_1 : boolean;
  signal LOAD_ncol_ind_611_load_0_req_0 : boolean;
  signal LOAD_ncol_ind_611_load_0_ack_0 : boolean;
  signal ptr_deref_816_load_0_ack_1 : boolean;
  signal LOAD_ncol_ind_611_load_0_req_1 : boolean;
  signal LOAD_ncol_ind_611_load_0_ack_1 : boolean;
  signal type_cast_615_inst_req_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal addr_of_812_final_reg_req_1 : boolean;
  signal ADD_u32_u32_620_inst_req_0 : boolean;
  signal ADD_u32_u32_620_inst_ack_0 : boolean;
  signal ADD_u32_u32_620_inst_req_1 : boolean;
  signal ADD_u32_u32_620_inst_ack_1 : boolean;
  signal ADD_u32_u32_626_inst_req_0 : boolean;
  signal ADD_u32_u32_626_inst_ack_0 : boolean;
  signal ADD_u32_u32_626_inst_req_1 : boolean;
  signal ADD_u32_u32_626_inst_ack_1 : boolean;
  signal SLT_i32_u1_633_inst_req_0 : boolean;
  signal SLT_i32_u1_633_inst_ack_0 : boolean;
  signal SLT_i32_u1_633_inst_req_1 : boolean;
  signal SLT_i32_u1_633_inst_ack_1 : boolean;
  signal addr_of_812_final_reg_req_0 : boolean;
  signal addr_of_812_final_reg_ack_0 : boolean;
  signal if_stmt_635_branch_req_0 : boolean;
  signal if_stmt_635_branch_ack_1 : boolean;
  signal if_stmt_635_branch_ack_0 : boolean;
  signal ptr_deref_644_load_0_req_0 : boolean;
  signal ptr_deref_644_load_0_ack_0 : boolean;
  signal ptr_deref_644_load_0_req_1 : boolean;
  signal ptr_deref_644_load_0_ack_1 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal type_cast_648_inst_req_1 : boolean;
  signal type_cast_648_inst_ack_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal addr_of_654_final_reg_req_0 : boolean;
  signal addr_of_654_final_reg_ack_0 : boolean;
  signal addr_of_654_final_reg_req_1 : boolean;
  signal addr_of_654_final_reg_ack_1 : boolean;
  signal ptr_deref_658_load_0_req_0 : boolean;
  signal ptr_deref_658_load_0_ack_0 : boolean;
  signal ptr_deref_658_load_0_req_1 : boolean;
  signal ptr_deref_658_load_0_ack_1 : boolean;
  signal ptr_deref_661_store_0_req_0 : boolean;
  signal ptr_deref_661_store_0_ack_0 : boolean;
  signal ptr_deref_666_load_0_req_1 : boolean;
  signal ptr_deref_666_load_0_ack_1 : boolean;
  signal WPIPE_mem_out_668_inst_req_0 : boolean;
  signal WPIPE_mem_out_668_inst_ack_0 : boolean;
  signal WPIPE_mem_out_668_inst_req_1 : boolean;
  signal WPIPE_mem_out_668_inst_ack_1 : boolean;
  signal ptr_deref_675_load_0_req_0 : boolean;
  signal ptr_deref_675_load_0_ack_0 : boolean;
  signal ptr_deref_675_load_0_req_1 : boolean;
  signal ptr_deref_675_load_0_ack_1 : boolean;
  signal ADD_u32_u32_681_inst_req_0 : boolean;
  signal ADD_u32_u32_681_inst_ack_0 : boolean;
  signal ADD_u32_u32_681_inst_req_1 : boolean;
  signal ADD_u32_u32_681_inst_ack_1 : boolean;
  signal ptr_deref_684_store_0_req_0 : boolean;
  signal ptr_deref_684_store_0_ack_0 : boolean;
  signal ptr_deref_684_store_0_req_1 : boolean;
  signal ptr_deref_684_store_0_ack_1 : boolean;
  signal ptr_deref_690_store_0_req_0 : boolean;
  signal ptr_deref_690_store_0_ack_0 : boolean;
  signal ptr_deref_690_store_0_req_1 : boolean;
  signal ptr_deref_690_store_0_ack_1 : boolean;
  signal ptr_deref_698_load_0_req_0 : boolean;
  signal ptr_deref_698_load_0_ack_0 : boolean;
  signal ptr_deref_698_load_0_req_1 : boolean;
  signal ptr_deref_698_load_0_ack_1 : boolean;
  signal LOAD_ncols_701_load_0_req_0 : boolean;
  signal LOAD_ncols_701_load_0_ack_0 : boolean;
  signal LOAD_ncols_701_load_0_req_1 : boolean;
  signal LOAD_ncols_701_load_0_ack_1 : boolean;
  signal type_cast_705_inst_req_0 : boolean;
  signal type_cast_705_inst_ack_0 : boolean;
  signal type_cast_705_inst_req_1 : boolean;
  signal type_cast_705_inst_ack_1 : boolean;
  signal SLT_i32_u1_712_inst_req_0 : boolean;
  signal SLT_i32_u1_712_inst_ack_0 : boolean;
  signal SLT_i32_u1_712_inst_req_1 : boolean;
  signal SLT_i32_u1_712_inst_ack_1 : boolean;
  signal if_stmt_714_branch_req_0 : boolean;
  signal if_stmt_714_branch_ack_1 : boolean;
  signal if_stmt_714_branch_ack_0 : boolean;
  signal ptr_deref_723_load_0_req_0 : boolean;
  signal ptr_deref_723_load_0_ack_0 : boolean;
  signal ptr_deref_723_load_0_req_1 : boolean;
  signal ptr_deref_723_load_0_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal type_cast_728_inst_req_0 : boolean;
  signal type_cast_728_inst_ack_0 : boolean;
  signal type_cast_728_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_1 : boolean;
  signal addr_of_733_final_reg_req_0 : boolean;
  signal addr_of_733_final_reg_ack_0 : boolean;
  signal addr_of_733_final_reg_req_1 : boolean;
  signal addr_of_733_final_reg_ack_1 : boolean;
  signal ptr_deref_737_load_0_req_0 : boolean;
  signal ptr_deref_737_load_0_ack_0 : boolean;
  signal ptr_deref_737_load_0_req_1 : boolean;
  signal ptr_deref_737_load_0_ack_1 : boolean;
  signal ptr_deref_740_store_0_req_0 : boolean;
  signal ptr_deref_740_store_0_ack_0 : boolean;
  signal ptr_deref_740_store_0_req_1 : boolean;
  signal ptr_deref_740_store_0_ack_1 : boolean;
  signal ptr_deref_745_load_0_req_0 : boolean;
  signal ptr_deref_745_load_0_ack_0 : boolean;
  signal ptr_deref_745_load_0_req_1 : boolean;
  signal ptr_deref_745_load_0_ack_1 : boolean;
  signal WPIPE_code_block_out_747_inst_req_0 : boolean;
  signal WPIPE_code_block_out_747_inst_ack_0 : boolean;
  signal WPIPE_code_block_out_747_inst_req_1 : boolean;
  signal WPIPE_code_block_out_747_inst_ack_1 : boolean;
  signal ptr_deref_754_load_0_req_0 : boolean;
  signal ptr_deref_754_load_0_ack_0 : boolean;
  signal ptr_deref_754_load_0_req_1 : boolean;
  signal ptr_deref_754_load_0_ack_1 : boolean;
  signal ADD_u32_u32_760_inst_req_0 : boolean;
  signal ADD_u32_u32_760_inst_ack_0 : boolean;
  signal ADD_u32_u32_760_inst_req_1 : boolean;
  signal ADD_u32_u32_760_inst_ack_1 : boolean;
  signal ptr_deref_816_load_0_ack_0 : boolean;
  signal ptr_deref_816_load_0_req_0 : boolean;
  signal ptr_deref_763_store_0_req_0 : boolean;
  signal ptr_deref_763_store_0_ack_0 : boolean;
  signal ptr_deref_763_store_0_req_1 : boolean;
  signal ptr_deref_763_store_0_ack_1 : boolean;
  signal addr_of_812_final_reg_ack_1 : boolean;
  signal ptr_deref_769_store_0_req_0 : boolean;
  signal ptr_deref_769_store_0_ack_0 : boolean;
  signal ptr_deref_769_store_0_req_1 : boolean;
  signal ptr_deref_769_store_0_ack_1 : boolean;
  signal ptr_deref_777_load_0_req_0 : boolean;
  signal ptr_deref_777_load_0_ack_0 : boolean;
  signal ptr_deref_777_load_0_req_1 : boolean;
  signal ptr_deref_777_load_0_ack_1 : boolean;
  signal LOAD_ncols_780_load_0_req_0 : boolean;
  signal LOAD_ncols_780_load_0_ack_0 : boolean;
  signal LOAD_ncols_780_load_0_req_1 : boolean;
  signal LOAD_ncols_780_load_0_ack_1 : boolean;
  signal type_cast_784_inst_req_0 : boolean;
  signal type_cast_784_inst_ack_0 : boolean;
  signal type_cast_784_inst_req_1 : boolean;
  signal type_cast_784_inst_ack_1 : boolean;
  signal SLT_i32_u1_791_inst_req_0 : boolean;
  signal SLT_i32_u1_791_inst_ack_0 : boolean;
  signal SLT_i32_u1_791_inst_req_1 : boolean;
  signal SLT_i32_u1_791_inst_ack_1 : boolean;
  signal if_stmt_793_branch_req_0 : boolean;
  signal if_stmt_793_branch_ack_1 : boolean;
  signal if_stmt_793_branch_ack_0 : boolean;
  signal ptr_deref_802_load_0_req_0 : boolean;
  signal ptr_deref_802_load_0_ack_0 : boolean;
  signal ptr_deref_802_load_0_req_1 : boolean;
  signal ptr_deref_802_load_0_ack_1 : boolean;
  signal type_cast_806_inst_req_0 : boolean;
  signal type_cast_806_inst_ack_0 : boolean;
  signal type_cast_806_inst_req_1 : boolean;
  signal type_cast_806_inst_ack_1 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal type_cast_807_inst_req_1 : boolean;
  signal type_cast_807_inst_ack_1 : boolean;
  signal ptr_deref_819_store_0_req_0 : boolean;
  signal ptr_deref_819_store_0_ack_0 : boolean;
  signal ptr_deref_819_store_0_req_1 : boolean;
  signal ptr_deref_819_store_0_ack_1 : boolean;
  signal ptr_deref_824_load_0_req_0 : boolean;
  signal ptr_deref_824_load_0_ack_0 : boolean;
  signal ptr_deref_824_load_0_req_1 : boolean;
  signal ptr_deref_824_load_0_ack_1 : boolean;
  signal WPIPE_aPriori_out_826_inst_req_0 : boolean;
  signal WPIPE_aPriori_out_826_inst_ack_0 : boolean;
  signal WPIPE_aPriori_out_826_inst_req_1 : boolean;
  signal WPIPE_aPriori_out_826_inst_ack_1 : boolean;
  signal ptr_deref_833_load_0_req_0 : boolean;
  signal ptr_deref_833_load_0_ack_0 : boolean;
  signal ptr_deref_833_load_0_req_1 : boolean;
  signal ptr_deref_833_load_0_ack_1 : boolean;
  signal ADD_u32_u32_839_inst_req_0 : boolean;
  signal ADD_u32_u32_839_inst_ack_0 : boolean;
  signal ADD_u32_u32_839_inst_req_1 : boolean;
  signal ADD_u32_u32_839_inst_ack_1 : boolean;
  signal ptr_deref_842_store_0_req_0 : boolean;
  signal ptr_deref_842_store_0_ack_0 : boolean;
  signal ptr_deref_842_store_0_req_1 : boolean;
  signal ptr_deref_842_store_0_ack_1 : boolean;
  signal ptr_deref_849_load_0_req_0 : boolean;
  signal ptr_deref_849_load_0_ack_0 : boolean;
  signal ptr_deref_849_load_0_req_1 : boolean;
  signal ptr_deref_849_load_0_ack_1 : boolean;
  signal memory_space_18_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_18_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_18_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_18_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_18_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_18_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_18_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_18_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_19_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_19_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_19_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_19_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_19_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_19_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_19_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_19_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_19_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_19_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_19_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_19_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_19_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_19_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_19_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_19_sc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_20_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_20_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_20_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_20_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_20_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_20_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_20_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_20_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_20_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_20_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_20_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_20_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_20_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_20_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_20_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_20_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_21_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_21_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_21_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_21_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_21_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_21_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_21_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_21_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_21_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_21_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_21_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_21_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_21_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_21_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_21_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_21_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_22_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_22_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_22_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_22_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_22_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_22_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_22_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_22_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_22_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_22_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_22_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_22_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_22_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_22_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_22_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_22_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "send_output_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  send_output_CP_3660_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "send_output_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= send_output_CP_3660_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= send_output_CP_3660_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= send_output_CP_3660_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  send_output_CP_3660: Block -- control-path 
    signal send_output_CP_3660_elements: BooleanArray(244 downto 0);
    -- 
  begin -- 
    send_output_CP_3660_elements(0) <= send_output_CP_3660_start;
    send_output_CP_3660_symbol <= send_output_CP_3660_elements(244);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_566/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	31 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596__entry__
      -- CP-element group 1: 	 branch_block_stmt_566/branch_block_stmt_566__entry__
      -- 
    send_output_CP_3660_elements(1) <= send_output_CP_3660_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	33 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	202 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_566/bb_0_bb_1
      -- CP-element group 2: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596__exit__
      -- 
    send_output_CP_3660_elements(2) <= send_output_CP_3660_elements(33);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	205 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	34 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634__entry__
      -- CP-element group 3: 	 branch_block_stmt_566/merge_stmt_598__exit__
      -- 
    send_output_CP_3660_elements(3) <= send_output_CP_3660_elements(205);
    -- CP-element group 4:  branch  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	52 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4: 	54 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_566/if_stmt_635__entry__
      -- CP-element group 4: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634__exit__
      -- 
    send_output_CP_3660_elements(4) <= send_output_CP_3660_elements(52);
    -- CP-element group 5:  merge  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	208 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	62 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667__entry__
      -- CP-element group 5: 	 branch_block_stmt_566/merge_stmt_641__exit__
      -- 
    send_output_CP_3660_elements(5) <= send_output_CP_3660_elements(208);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	80 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	81 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_566/assign_stmt_670__entry__
      -- CP-element group 6: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667__exit__
      -- 
    send_output_CP_3660_elements(6) <= send_output_CP_3660_elements(80);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	83 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	209 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_566/bb_2_bb_3
      -- CP-element group 7: 	 branch_block_stmt_566/assign_stmt_670__exit__
      -- 
    send_output_CP_3660_elements(7) <= send_output_CP_3660_elements(83);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	211 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	84 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686__entry__
      -- CP-element group 8: 	 branch_block_stmt_566/merge_stmt_672__exit__
      -- 
    send_output_CP_3660_elements(8) <= send_output_CP_3660_elements(211);
    -- CP-element group 9:  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	91 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	203 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686__exit__
      -- CP-element group 9: 	 branch_block_stmt_566/bb_3_bb_1
      -- 
    send_output_CP_3660_elements(9) <= send_output_CP_3660_elements(91);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	214 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	93 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_566/merge_stmt_688__exit__
      -- CP-element group 10: 	 branch_block_stmt_566/assign_stmt_693__entry__
      -- 
    send_output_CP_3660_elements(10) <= send_output_CP_3660_elements(214);
    -- CP-element group 11:  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	95 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	215 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_566/bb_4_bb_5
      -- CP-element group 11: 	 branch_block_stmt_566/assign_stmt_693__exit__
      -- 
    send_output_CP_3660_elements(11) <= send_output_CP_3660_elements(95);
    -- CP-element group 12:  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	218 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713__entry__
      -- CP-element group 12: 	 branch_block_stmt_566/merge_stmt_695__exit__
      -- 
    send_output_CP_3660_elements(12) <= send_output_CP_3660_elements(218);
    -- CP-element group 13:  branch  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	105 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	106 
    -- CP-element group 13: 	107 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713__exit__
      -- CP-element group 13: 	 branch_block_stmt_566/if_stmt_714__entry__
      -- 
    send_output_CP_3660_elements(13) <= send_output_CP_3660_elements(105);
    -- CP-element group 14:  merge  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	221 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	115 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_566/merge_stmt_720__exit__
      -- CP-element group 14: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746__entry__
      -- 
    send_output_CP_3660_elements(14) <= send_output_CP_3660_elements(221);
    -- CP-element group 15:  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	133 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	134 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746__exit__
      -- CP-element group 15: 	 branch_block_stmt_566/assign_stmt_749__entry__
      -- 
    send_output_CP_3660_elements(15) <= send_output_CP_3660_elements(133);
    -- CP-element group 16:  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	136 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	222 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_566/bb_6_bb_7
      -- CP-element group 16: 	 branch_block_stmt_566/assign_stmt_749__exit__
      -- 
    send_output_CP_3660_elements(16) <= send_output_CP_3660_elements(136);
    -- CP-element group 17:  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	224 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	137 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765__entry__
      -- CP-element group 17: 	 branch_block_stmt_566/merge_stmt_751__exit__
      -- 
    send_output_CP_3660_elements(17) <= send_output_CP_3660_elements(224);
    -- CP-element group 18:  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	144 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	216 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_566/bb_7_bb_5
      -- CP-element group 18: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765__exit__
      -- 
    send_output_CP_3660_elements(18) <= send_output_CP_3660_elements(144);
    -- CP-element group 19:  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	227 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	146 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_566/assign_stmt_772__entry__
      -- CP-element group 19: 	 branch_block_stmt_566/merge_stmt_767__exit__
      -- 
    send_output_CP_3660_elements(19) <= send_output_CP_3660_elements(227);
    -- CP-element group 20:  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	148 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	229 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_566/bb_8_bb_9
      -- CP-element group 20: 	 branch_block_stmt_566/assign_stmt_772__exit__
      -- 
    send_output_CP_3660_elements(20) <= send_output_CP_3660_elements(148);
    -- CP-element group 21:  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	231 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	149 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792__entry__
      -- CP-element group 21: 	 branch_block_stmt_566/merge_stmt_774__exit__
      -- 
    send_output_CP_3660_elements(21) <= send_output_CP_3660_elements(231);
    -- CP-element group 22:  branch  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	158 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	159 
    -- CP-element group 22: 	160 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_566/if_stmt_793__entry__
      -- CP-element group 22: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792__exit__
      -- 
    send_output_CP_3660_elements(22) <= send_output_CP_3660_elements(158);
    -- CP-element group 23:  merge  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	234 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	168 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825__entry__
      -- CP-element group 23: 	 branch_block_stmt_566/merge_stmt_799__exit__
      -- 
    send_output_CP_3660_elements(23) <= send_output_CP_3660_elements(234);
    -- CP-element group 24:  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	186 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	187 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_566/assign_stmt_828__entry__
      -- CP-element group 24: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825__exit__
      -- 
    send_output_CP_3660_elements(24) <= send_output_CP_3660_elements(186);
    -- CP-element group 25:  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	189 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	235 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_566/bb_10_bb_11
      -- CP-element group 25: 	 branch_block_stmt_566/assign_stmt_828__exit__
      -- 
    send_output_CP_3660_elements(25) <= send_output_CP_3660_elements(189);
    -- CP-element group 26:  place  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	237 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	190 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_566/merge_stmt_830__exit__
      -- CP-element group 26: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844__entry__
      -- 
    send_output_CP_3660_elements(26) <= send_output_CP_3660_elements(237);
    -- CP-element group 27:  place  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	197 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	228 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_566/bb_11_bb_9
      -- CP-element group 27: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844__exit__
      -- 
    send_output_CP_3660_elements(27) <= send_output_CP_3660_elements(197);
    -- CP-element group 28:  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	240 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	199 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_566/merge_stmt_846__exit__
      -- CP-element group 28: 	 branch_block_stmt_566/assign_stmt_850__entry__
      -- 
    send_output_CP_3660_elements(28) <= send_output_CP_3660_elements(240);
    -- CP-element group 29:  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	201 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	241 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_566/assign_stmt_850__exit__
      -- CP-element group 29: 	 branch_block_stmt_566/return__
      -- 
    send_output_CP_3660_elements(29) <= send_output_CP_3660_elements(201);
    -- CP-element group 30:  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	243 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	244 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_566/merge_stmt_852__exit__
      -- CP-element group 30: 	 branch_block_stmt_566/branch_block_stmt_566__exit__
      -- 
    send_output_CP_3660_elements(30) <= send_output_CP_3660_elements(243);
    -- CP-element group 31:  fork  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (31) 
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_word_addrgen/$exit
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_update_start_
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/ptr_deref_593_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/ptr_deref_593_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/word_0/cr
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_word_addrgen/root_register_req
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/ptr_deref_593_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/ptr_deref_593_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_addr_resize/base_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_addr_resize/base_resize_req
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_addr_resize/$exit
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_addr_resize/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_word_addrgen/root_register_ack
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_base_address_resized
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_word_addrgen/$entry
      -- 
    cr_3783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(31), ack => ptr_deref_593_store_0_req_1); -- 
    rr_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(31), ack => ptr_deref_593_store_0_req_0); -- 
    send_output_CP_3660_elements(31) <= send_output_CP_3660_elements(1);
    -- CP-element group 32:  transition  input  no-bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Sample/word_access_start/word_0/ra
      -- 
    ra_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_store_0_ack_0, ack => send_output_CP_3660_elements(32)); -- 
    -- CP-element group 33:  transition  input  no-bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	2 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/$exit
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/word_0/ca
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_566/assign_stmt_575_to_assign_stmt_596/ptr_deref_593_Update/word_access_complete/word_0/$exit
      -- 
    ca_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_store_0_ack_1, ack => send_output_CP_3660_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	3 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34: 	44 
    -- CP-element group 34: 	47 
    -- CP-element group 34: 	49 
    -- CP-element group 34: 	52 
    -- CP-element group 34:  members (66) 
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_word_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_root_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_address_resized
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_addr_resize/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_addr_resize/$exit
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_addr_resize/base_resize_req
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_addr_resize/base_resize_ack
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_plus_offset/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_plus_offset/$exit
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_plus_offset/sum_rename_req
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_base_plus_offset/sum_rename_ack
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_word_addrgen/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_word_addrgen/$exit
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_word_addrgen/root_register_req
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_word_addrgen/root_register_ack
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/word_0/rr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/word_0/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_word_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_root_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/word_0/rr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/word_0/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_word_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_root_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/word_0/rr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/word_0/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_update_start_
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Update/cr
      -- 
    cr_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => ptr_deref_601_load_0_req_1); -- 
    rr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => ptr_deref_601_load_0_req_0); -- 
    cr_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => LOAD_nrows_604_load_0_req_1); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => LOAD_nrows_604_load_0_req_0); -- 
    cr_3883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => type_cast_608_inst_req_1); -- 
    cr_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => LOAD_ncol_ind_611_load_0_req_1); -- 
    rr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => LOAD_ncol_ind_611_load_0_req_0); -- 
    cr_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => type_cast_615_inst_req_1); -- 
    cr_3944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => ADD_u32_u32_620_inst_req_1); -- 
    cr_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => ADD_u32_u32_626_inst_req_1); -- 
    cr_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(34), ack => SLT_i32_u1_633_inst_req_1); -- 
    send_output_CP_3660_elements(34) <= send_output_CP_3660_elements(3);
    -- CP-element group 35:  transition  input  no-bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Sample/word_access_start/word_0/ra
      -- 
    ra_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_601_load_0_ack_0, ack => send_output_CP_3660_elements(35)); -- 
    -- CP-element group 36:  transition  input  no-bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	50 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/word_access_complete/word_0/ca
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/ptr_deref_601_Merge/$entry
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/ptr_deref_601_Merge/$exit
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/ptr_deref_601_Merge/merge_req
      -- CP-element group 36: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ptr_deref_601_Update/ptr_deref_601_Merge/merge_ack
      -- 
    ca_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_601_load_0_ack_1, ack => send_output_CP_3660_elements(36)); -- 
    -- CP-element group 37:  transition  input  no-bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/$exit
      -- CP-element group 37: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Sample/word_access_start/word_0/ra
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_604_load_0_ack_0, ack => send_output_CP_3660_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  no-bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (12) 
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/word_access_complete/word_0/ca
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/LOAD_nrows_604_Merge/$entry
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/LOAD_nrows_604_Merge/$exit
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/LOAD_nrows_604_Merge/merge_req
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_nrows_604_Update/LOAD_nrows_604_Merge/merge_ack
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Sample/rr
      -- 
    ca_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_604_load_0_ack_1, ack => send_output_CP_3660_elements(38)); -- 
    rr_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(38), ack => type_cast_608_inst_req_0); -- 
    -- CP-element group 39:  transition  input  no-bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Sample/ra
      -- 
    ra_3879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => send_output_CP_3660_elements(39)); -- 
    -- CP-element group 40:  transition  input  no-bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	45 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_608_Update/ca
      -- 
    ca_3884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => send_output_CP_3660_elements(40)); -- 
    -- CP-element group 41:  transition  input  no-bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/$exit
      -- CP-element group 41: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Sample/word_access_start/word_0/ra
      -- 
    ra_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_611_load_0_ack_0, ack => send_output_CP_3660_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  no-bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (12) 
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/word_access_complete/word_0/ca
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/LOAD_ncol_ind_611_Merge/$entry
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/LOAD_ncol_ind_611_Merge/$exit
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/LOAD_ncol_ind_611_Merge/merge_req
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/LOAD_ncol_ind_611_Update/LOAD_ncol_ind_611_Merge/merge_ack
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Sample/rr
      -- 
    ca_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_611_load_0_ack_1, ack => send_output_CP_3660_elements(42)); -- 
    rr_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(42), ack => type_cast_615_inst_req_0); -- 
    -- CP-element group 43:  transition  input  no-bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Sample/ra
      -- 
    ra_3926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => send_output_CP_3660_elements(43)); -- 
    -- CP-element group 44:  transition  input  no-bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	34 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/type_cast_615_Update/ca
      -- 
    ca_3931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => send_output_CP_3660_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	40 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Sample/rr
      -- 
    rr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(45), ack => ADD_u32_u32_620_inst_req_0); -- 
    send_output_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(40) & send_output_CP_3660_elements(44);
      gj_send_output_cp_element_group_45 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  no-bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Sample/ra
      -- 
    ra_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_620_inst_ack_0, ack => send_output_CP_3660_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  no-bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	34 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_620_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Sample/rr
      -- 
    ca_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_620_inst_ack_1, ack => send_output_CP_3660_elements(47)); -- 
    rr_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(47), ack => ADD_u32_u32_626_inst_req_0); -- 
    -- CP-element group 48:  transition  input  no-bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Sample/ra
      -- 
    ra_3954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_626_inst_ack_0, ack => send_output_CP_3660_elements(48)); -- 
    -- CP-element group 49:  transition  input  no-bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	34 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/ADD_u32_u32_626_Update/ca
      -- 
    ca_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_626_inst_ack_1, ack => send_output_CP_3660_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	36 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Sample/rr
      -- 
    rr_3967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(50), ack => SLT_i32_u1_633_inst_req_0); -- 
    send_output_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(36) & send_output_CP_3660_elements(49);
      gj_send_output_cp_element_group_50 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  no-bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Sample/ra
      -- 
    ra_3968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_633_inst_ack_0, ack => send_output_CP_3660_elements(51)); -- 
    -- CP-element group 52:  transition  input  no-bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	34 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	4 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/$exit
      -- CP-element group 52: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_566/assign_stmt_602_to_assign_stmt_634/SLT_i32_u1_633_Update/ca
      -- 
    ca_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_633_inst_ack_1, ack => send_output_CP_3660_elements(52)); -- 
    -- CP-element group 53:  transition  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_566/if_stmt_635_dead_link/$entry
      -- 
    send_output_CP_3660_elements(53) <= send_output_CP_3660_elements(4);
    -- CP-element group 54:  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	4 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_566/if_stmt_635_eval_test/$entry
      -- CP-element group 54: 	 branch_block_stmt_566/if_stmt_635_eval_test/$exit
      -- CP-element group 54: 	 branch_block_stmt_566/if_stmt_635_eval_test/branch_req
      -- 
    branch_req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(54), ack => if_stmt_635_branch_req_0); -- 
    send_output_CP_3660_elements(54) <= send_output_CP_3660_elements(4);
    -- CP-element group 55:  branch  place  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_566/R_iNsTr_10_636_place
      -- 
    send_output_CP_3660_elements(55) <= send_output_CP_3660_elements(54);
    -- CP-element group 56:  transition  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_566/if_stmt_635_if_link/$entry
      -- 
    send_output_CP_3660_elements(56) <= send_output_CP_3660_elements(55);
    -- CP-element group 57:  transition  input  no-bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_566/if_stmt_635_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_566/if_stmt_635_if_link/if_choice_transition
      -- 
    if_choice_transition_3986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_635_branch_ack_1, ack => send_output_CP_3660_elements(57)); -- 
    -- CP-element group 58:  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_566/if_stmt_635_else_link/$entry
      -- 
    send_output_CP_3660_elements(58) <= send_output_CP_3660_elements(55);
    -- CP-element group 59:  transition  input  no-bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_566/if_stmt_635_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_566/if_stmt_635_else_link/else_choice_transition
      -- 
    else_choice_transition_3990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_635_branch_ack_0, ack => send_output_CP_3660_elements(59)); -- 
    -- CP-element group 60:  place  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	57 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	206 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_566/bb_1_bb_2
      -- 
    send_output_CP_3660_elements(60) <= send_output_CP_3660_elements(57);
    -- CP-element group 61:  place  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	212 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_566/bb_1_bb_4
      -- 
    send_output_CP_3660_elements(61) <= send_output_CP_3660_elements(59);
    -- CP-element group 62:  join  fork  transition  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	5 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	68 
    -- CP-element group 62: 	70 
    -- CP-element group 62: 	72 
    -- CP-element group 62: 	73 
    -- CP-element group 62: 	75 
    -- CP-element group 62: 	76 
    -- CP-element group 62: 	78 
    -- CP-element group 62:  members (83) 
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/word_0/rr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_complete/req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_update_start_
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/word_0/cr
      -- 
    cr_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => ptr_deref_644_load_0_req_1); -- 
    rr_4028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => ptr_deref_644_load_0_req_0); -- 
    cr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => type_cast_649_inst_req_1); -- 
    cr_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => type_cast_648_inst_req_1); -- 
    req_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => addr_of_654_final_reg_req_1); -- 
    cr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => ptr_deref_658_load_0_req_1); -- 
    cr_4211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => ptr_deref_661_store_0_req_1); -- 
    cr_4256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(62), ack => ptr_deref_666_load_0_req_1); -- 
    send_output_CP_3660_elements(62) <= send_output_CP_3660_elements(5);
    -- CP-element group 63:  transition  input  no-bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Sample/word_access_start/word_0/ra
      -- 
    ra_4029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_load_0_ack_0, ack => send_output_CP_3660_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  no-bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (12) 
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/ptr_deref_644_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/ptr_deref_644_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/ptr_deref_644_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_644_Update/ptr_deref_644_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Sample/rr
      -- 
    ca_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_load_0_ack_1, ack => send_output_CP_3660_elements(64)); -- 
    rr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(64), ack => type_cast_648_inst_req_0); -- 
    -- CP-element group 65:  transition  input  no-bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Sample/ra
      -- 
    ra_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_0, ack => send_output_CP_3660_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  no-bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_648_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Sample/rr
      -- 
    ca_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_1, ack => send_output_CP_3660_elements(66)); -- 
    rr_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(66), ack => type_cast_649_inst_req_0); -- 
    -- CP-element group 67:  transition  input  no-bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Sample/ra
      -- 
    ra_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => send_output_CP_3660_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  no-bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	62 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (27) 
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/type_cast_649_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_resized_0
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_scaled_0
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_computed_0
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_resize_0/$entry
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_resize_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_resize_0/index_resize_req
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_resize_0/index_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_scale_0/$entry
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_scale_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_scale_0/scale_rename_req
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_index_scale_0/scale_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_final_index_sum_regn/$entry
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_final_index_sum_regn/$exit
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_final_index_sum_regn/req
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_final_index_sum_regn/ack
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/array_obj_ref_653_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_request/req
      -- 
    ca_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => send_output_CP_3660_elements(68)); -- 
    req_4106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(68), ack => addr_of_654_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  no-bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	80 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_request/ack
      -- 
    ack_4107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_0, ack => send_output_CP_3660_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	62 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (24) 
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/addr_of_654_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_word_addrgen/root_register_ack
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/word_0/$entry
      -- CP-element group 70: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/word_0/rr
      -- 
    ack_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_1, ack => send_output_CP_3660_elements(70)); -- 
    rr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(70), ack => ptr_deref_658_load_0_req_0); -- 
    -- CP-element group 71:  transition  input  no-bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/$exit
      -- CP-element group 71: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Sample/word_access_start/word_0/ra
      -- 
    ra_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_load_0_ack_0, ack => send_output_CP_3660_elements(71)); -- 
    -- CP-element group 72:  transition  input  no-bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	62 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (9) 
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/word_access_complete/word_0/ca
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/ptr_deref_658_Merge/$entry
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/ptr_deref_658_Merge/$exit
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/ptr_deref_658_Merge/merge_req
      -- CP-element group 72: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_658_Update/ptr_deref_658_Merge/merge_ack
      -- 
    ca_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_load_0_ack_1, ack => send_output_CP_3660_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  no-bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	62 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/ptr_deref_661_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/ptr_deref_661_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/ptr_deref_661_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/ptr_deref_661_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/word_0/rr
      -- 
    rr_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(73), ack => ptr_deref_661_store_0_req_0); -- 
    send_output_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(62) & send_output_CP_3660_elements(72);
      gj_send_output_cp_element_group_73 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  no-bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	79 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Sample/word_access_start/word_0/ra
      -- 
    ra_4201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_store_0_ack_0, ack => send_output_CP_3660_elements(74)); -- 
    -- CP-element group 75:  transition  input  no-bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	62 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/word_0/ca
      -- CP-element group 75: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_update_completed_
      -- 
    ca_4212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_store_0_ack_1, ack => send_output_CP_3660_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  no-bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	62 
    -- CP-element group 76: 	79 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/word_0/rr
      -- CP-element group 76: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/$entry
      -- CP-element group 76: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_sample_start_
      -- 
    rr_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(76), ack => ptr_deref_666_load_0_req_0); -- 
    send_output_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(62) & send_output_CP_3660_elements(79);
      gj_send_output_cp_element_group_76 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  no-bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/$exit
      -- CP-element group 77: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/word_access_start/word_0/ra
      -- CP-element group 77: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Sample/$exit
      -- 
    ra_4246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_666_load_0_ack_0, ack => send_output_CP_3660_elements(77)); -- 
    -- CP-element group 78:  transition  input  no-bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	62 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/$exit
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/word_access_complete/word_0/ca
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/ptr_deref_666_Merge/$entry
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/ptr_deref_666_Merge/$exit
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/ptr_deref_666_Merge/merge_req
      -- CP-element group 78: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_666_Update/ptr_deref_666_Merge/merge_ack
      -- 
    ca_4257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_666_load_0_ack_1, ack => send_output_CP_3660_elements(78)); -- 
    -- CP-element group 79:  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	76 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/ptr_deref_661_ptr_deref_666_delay
      -- 
    -- Element group send_output_CP_3660_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(74), ack => send_output_CP_3660_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  transition  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	69 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	6 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_566/assign_stmt_645_to_assign_stmt_667/$exit
      -- 
    send_output_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(69) & send_output_CP_3660_elements(75) & send_output_CP_3660_elements(78);
      gj_send_output_cp_element_group_80 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	6 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_566/assign_stmt_670/$entry
      -- CP-element group 81: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Sample/req
      -- 
    req_4274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(81), ack => WPIPE_mem_out_668_inst_req_0); -- 
    send_output_CP_3660_elements(81) <= send_output_CP_3660_elements(6);
    -- CP-element group 82:  transition  input  output  no-bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_update_start_
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Sample/ack
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Update/req
      -- 
    ack_4275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_out_668_inst_ack_0, ack => send_output_CP_3660_elements(82)); -- 
    req_4279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(82), ack => WPIPE_mem_out_668_inst_req_1); -- 
    -- CP-element group 83:  transition  input  no-bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	7 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_566/assign_stmt_670/$exit
      -- CP-element group 83: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_566/assign_stmt_670/WPIPE_mem_out_668_Update/ack
      -- 
    ack_4280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_out_668_inst_ack_1, ack => send_output_CP_3660_elements(83)); -- 
    -- CP-element group 84:  join  fork  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84: 	88 
    -- CP-element group 84: 	89 
    -- CP-element group 84: 	91 
    -- CP-element group 84:  members (51) 
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_update_start_
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_word_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_root_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_address_resized
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_addr_resize/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_addr_resize/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_addr_resize/base_resize_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_addr_resize/base_resize_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_plus_offset/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_plus_offset/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_plus_offset/sum_rename_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_base_plus_offset/sum_rename_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_word_addrgen/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_word_addrgen/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_word_addrgen/root_register_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_word_addrgen/root_register_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/word_0/rr
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/word_0/cr
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_update_start_
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Update/cr
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_update_start_
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_word_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_root_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_address_resized
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_addr_resize/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_addr_resize/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_addr_resize/base_resize_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_addr_resize/base_resize_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_plus_offset/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_plus_offset/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_plus_offset/sum_rename_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_base_plus_offset/sum_rename_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_word_addrgen/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_word_addrgen/$exit
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_word_addrgen/root_register_req
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_word_addrgen/root_register_ack
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/word_0/cr
      -- 
    cr_4327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(84), ack => ptr_deref_675_load_0_req_1); -- 
    rr_4316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(84), ack => ptr_deref_675_load_0_req_0); -- 
    cr_4346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(84), ack => ADD_u32_u32_681_inst_req_1); -- 
    cr_4396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(84), ack => ptr_deref_684_store_0_req_1); -- 
    send_output_CP_3660_elements(84) <= send_output_CP_3660_elements(8);
    -- CP-element group 85:  transition  input  no-bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	92 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/$exit
      -- CP-element group 85: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Sample/word_access_start/word_0/ra
      -- 
    ra_4317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_675_load_0_ack_0, ack => send_output_CP_3660_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  no-bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (12) 
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/word_access_complete/word_0/ca
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/ptr_deref_675_Merge/$entry
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/ptr_deref_675_Merge/$exit
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/ptr_deref_675_Merge/merge_req
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_Update/ptr_deref_675_Merge/merge_ack
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Sample/rr
      -- 
    ca_4328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_675_load_0_ack_1, ack => send_output_CP_3660_elements(86)); -- 
    rr_4341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(86), ack => ADD_u32_u32_681_inst_req_0); -- 
    -- CP-element group 87:  transition  input  no-bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Sample/ra
      -- 
    ra_4342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_681_inst_ack_0, ack => send_output_CP_3660_elements(87)); -- 
    -- CP-element group 88:  transition  input  no-bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ADD_u32_u32_681_Update/ca
      -- 
    ca_4347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_681_inst_ack_1, ack => send_output_CP_3660_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  no-bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	84 
    -- CP-element group 89: 	88 
    -- CP-element group 89: 	92 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/ptr_deref_684_Split/$entry
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/ptr_deref_684_Split/$exit
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/ptr_deref_684_Split/split_req
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/ptr_deref_684_Split/split_ack
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/word_0/rr
      -- 
    rr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(89), ack => ptr_deref_684_store_0_req_0); -- 
    send_output_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 31) := "send_output_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(84) & send_output_CP_3660_elements(88) & send_output_CP_3660_elements(92);
      gj_send_output_cp_element_group_89 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  no-bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/$exit
      -- CP-element group 90: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Sample/word_access_start/word_0/ra
      -- 
    ra_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_684_store_0_ack_0, ack => send_output_CP_3660_elements(90)); -- 
    -- CP-element group 91:  transition  input  no-bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	84 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	9 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/$exit
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/$exit
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_684_Update/word_access_complete/word_0/ca
      -- 
    ca_4397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_684_store_0_ack_1, ack => send_output_CP_3660_elements(91)); -- 
    -- CP-element group 92:  transition  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	85 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	89 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_566/assign_stmt_676_to_assign_stmt_686/ptr_deref_675_ptr_deref_684_delay
      -- 
    -- Element group send_output_CP_3660_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(85), ack => send_output_CP_3660_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	10 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (31) 
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_update_start_
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_address_calculated
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_word_address_calculated
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_root_address_calculated
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_address_resized
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_addr_resize/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_addr_resize/$exit
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_addr_resize/base_resize_req
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_addr_resize/base_resize_ack
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_plus_offset/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_plus_offset/$exit
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_plus_offset/sum_rename_req
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_base_plus_offset/sum_rename_ack
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_word_addrgen/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_word_addrgen/$exit
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_word_addrgen/root_register_req
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_word_addrgen/root_register_ack
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/ptr_deref_690_Split/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/ptr_deref_690_Split/$exit
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/ptr_deref_690_Split/split_req
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/ptr_deref_690_Split/split_ack
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/word_0/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/word_0/rr
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/word_0/$entry
      -- CP-element group 93: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/word_0/cr
      -- 
    cr_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(93), ack => ptr_deref_690_store_0_req_1); -- 
    rr_4439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(93), ack => ptr_deref_690_store_0_req_0); -- 
    send_output_CP_3660_elements(93) <= send_output_CP_3660_elements(10);
    -- CP-element group 94:  transition  input  no-bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/$exit
      -- CP-element group 94: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Sample/word_access_start/word_0/ra
      -- 
    ra_4440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_690_store_0_ack_0, ack => send_output_CP_3660_elements(94)); -- 
    -- CP-element group 95:  transition  input  no-bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	11 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/$exit
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/$exit
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_566/assign_stmt_693/ptr_deref_690_Update/word_access_complete/word_0/ca
      -- 
    ca_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_690_store_0_ack_1, ack => send_output_CP_3660_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	98 
    -- CP-element group 96: 	99 
    -- CP-element group 96: 	100 
    -- CP-element group 96: 	102 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (45) 
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_update_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_word_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_root_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_address_resized
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_addr_resize/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_addr_resize/$exit
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_addr_resize/base_resize_req
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_addr_resize/base_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_plus_offset/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_plus_offset/$exit
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_plus_offset/sum_rename_req
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_base_plus_offset/sum_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_word_addrgen/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_word_addrgen/$exit
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_word_addrgen/root_register_req
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_word_addrgen/root_register_ack
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/word_0/rr
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/word_0/cr
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_update_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_word_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_root_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/word_0/rr
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/word_0/cr
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_update_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Update/cr
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_update_start_
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Update/cr
      -- 
    cr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => ptr_deref_698_load_0_req_1); -- 
    rr_4487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => ptr_deref_698_load_0_req_0); -- 
    cr_4531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => LOAD_ncols_701_load_0_req_1); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => LOAD_ncols_701_load_0_req_0); -- 
    cr_4550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => type_cast_705_inst_req_1); -- 
    cr_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(96), ack => SLT_i32_u1_712_inst_req_1); -- 
    send_output_CP_3660_elements(96) <= send_output_CP_3660_elements(12);
    -- CP-element group 97:  transition  input  no-bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Sample/word_access_start/word_0/ra
      -- 
    ra_4488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_698_load_0_ack_0, ack => send_output_CP_3660_elements(97)); -- 
    -- CP-element group 98:  transition  input  no-bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/ptr_deref_698_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/ptr_deref_698_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/ptr_deref_698_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/ptr_deref_698_Update/ptr_deref_698_Merge/merge_ack
      -- 
    ca_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_698_load_0_ack_1, ack => send_output_CP_3660_elements(98)); -- 
    -- CP-element group 99:  transition  input  no-bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Sample/word_access_start/word_0/ra
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_701_load_0_ack_0, ack => send_output_CP_3660_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  no-bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (12) 
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/LOAD_ncols_701_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/LOAD_ncols_701_Merge/$exit
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/LOAD_ncols_701_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/LOAD_ncols_701_Update/LOAD_ncols_701_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Sample/rr
      -- 
    ca_4532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_701_load_0_ack_1, ack => send_output_CP_3660_elements(100)); -- 
    rr_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(100), ack => type_cast_705_inst_req_0); -- 
    -- CP-element group 101:  transition  input  no-bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Sample/ra
      -- 
    ra_4546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_0, ack => send_output_CP_3660_elements(101)); -- 
    -- CP-element group 102:  transition  input  no-bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	96 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/type_cast_705_Update/ca
      -- 
    ca_4551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_1, ack => send_output_CP_3660_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Sample/rr
      -- 
    rr_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(103), ack => SLT_i32_u1_712_inst_req_0); -- 
    send_output_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(98) & send_output_CP_3660_elements(102);
      gj_send_output_cp_element_group_103 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  no-bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Sample/ra
      -- 
    ra_4560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_712_inst_ack_0, ack => send_output_CP_3660_elements(104)); -- 
    -- CP-element group 105:  transition  input  no-bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	13 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/$exit
      -- CP-element group 105: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_566/assign_stmt_699_to_assign_stmt_713/SLT_i32_u1_712_Update/ca
      -- 
    ca_4565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_712_inst_ack_1, ack => send_output_CP_3660_elements(105)); -- 
    -- CP-element group 106:  transition  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	13 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_566/if_stmt_714_dead_link/$entry
      -- 
    send_output_CP_3660_elements(106) <= send_output_CP_3660_elements(13);
    -- CP-element group 107:  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	13 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_566/if_stmt_714_eval_test/$entry
      -- CP-element group 107: 	 branch_block_stmt_566/if_stmt_714_eval_test/$exit
      -- CP-element group 107: 	 branch_block_stmt_566/if_stmt_714_eval_test/branch_req
      -- 
    branch_req_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(107), ack => if_stmt_714_branch_req_0); -- 
    send_output_CP_3660_elements(107) <= send_output_CP_3660_elements(13);
    -- CP-element group 108:  branch  place  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_566/R_iNsTr_31_715_place
      -- 
    send_output_CP_3660_elements(108) <= send_output_CP_3660_elements(107);
    -- CP-element group 109:  transition  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_566/if_stmt_714_if_link/$entry
      -- 
    send_output_CP_3660_elements(109) <= send_output_CP_3660_elements(108);
    -- CP-element group 110:  transition  input  no-bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_566/if_stmt_714_if_link/$exit
      -- CP-element group 110: 	 branch_block_stmt_566/if_stmt_714_if_link/if_choice_transition
      -- 
    if_choice_transition_4578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_714_branch_ack_1, ack => send_output_CP_3660_elements(110)); -- 
    -- CP-element group 111:  transition  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_566/if_stmt_714_else_link/$entry
      -- 
    send_output_CP_3660_elements(111) <= send_output_CP_3660_elements(108);
    -- CP-element group 112:  transition  input  no-bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_566/if_stmt_714_else_link/$exit
      -- CP-element group 112: 	 branch_block_stmt_566/if_stmt_714_else_link/else_choice_transition
      -- 
    else_choice_transition_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_714_branch_ack_0, ack => send_output_CP_3660_elements(112)); -- 
    -- CP-element group 113:  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	219 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_566/bb_5_bb_6
      -- 
    send_output_CP_3660_elements(113) <= send_output_CP_3660_elements(110);
    -- CP-element group 114:  place  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	225 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_566/bb_5_bb_8
      -- 
    send_output_CP_3660_elements(114) <= send_output_CP_3660_elements(112);
    -- CP-element group 115:  join  fork  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	117 
    -- CP-element group 115: 	119 
    -- CP-element group 115: 	121 
    -- CP-element group 115: 	123 
    -- CP-element group 115: 	125 
    -- CP-element group 115: 	126 
    -- CP-element group 115: 	128 
    -- CP-element group 115: 	129 
    -- CP-element group 115: 	131 
    -- CP-element group 115:  members (83) 
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_word_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_root_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_address_resized
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_addr_resize/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_addr_resize/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_addr_resize/base_resize_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_addr_resize/base_resize_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_plus_offset/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_plus_offset/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_plus_offset/sum_rename_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_base_plus_offset/sum_rename_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_word_addrgen/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_word_addrgen/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_word_addrgen/root_register_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_word_addrgen/root_register_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/word_0/rr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/word_0/cr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_complete/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_complete/req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/word_0/cr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_word_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_root_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_address_resized
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_addr_resize/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_addr_resize/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_addr_resize/base_resize_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_addr_resize/base_resize_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_plus_offset/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_plus_offset/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_plus_offset/sum_rename_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_base_plus_offset/sum_rename_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_word_addrgen/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_word_addrgen/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_word_addrgen/root_register_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_word_addrgen/root_register_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/word_0/cr
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_update_start_
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_word_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_root_address_calculated
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_address_resized
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_addr_resize/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_addr_resize/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_addr_resize/base_resize_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_addr_resize/base_resize_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_plus_offset/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_plus_offset/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_plus_offset/sum_rename_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_base_plus_offset/sum_rename_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_word_addrgen/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_word_addrgen/$exit
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_word_addrgen/root_register_req
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_word_addrgen/root_register_ack
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/word_0/cr
      -- 
    cr_4631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => ptr_deref_723_load_0_req_1); -- 
    rr_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => ptr_deref_723_load_0_req_0); -- 
    cr_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => type_cast_728_inst_req_1); -- 
    cr_4654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => type_cast_727_inst_req_1); -- 
    req_4703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => addr_of_733_final_reg_req_1); -- 
    cr_4748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => ptr_deref_737_load_0_req_1); -- 
    cr_4803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => ptr_deref_740_store_0_req_1); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(115), ack => ptr_deref_745_load_0_req_1); -- 
    send_output_CP_3660_elements(115) <= send_output_CP_3660_elements(14);
    -- CP-element group 116:  transition  input  no-bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/$exit
      -- CP-element group 116: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Sample/word_access_start/word_0/ra
      -- 
    ra_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_723_load_0_ack_0, ack => send_output_CP_3660_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  no-bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (12) 
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/$exit
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/word_access_complete/word_0/ca
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/ptr_deref_723_Merge/$entry
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/ptr_deref_723_Merge/$exit
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/ptr_deref_723_Merge/merge_req
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_723_Update/ptr_deref_723_Merge/merge_ack
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Sample/rr
      -- 
    ca_4632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_723_load_0_ack_1, ack => send_output_CP_3660_elements(117)); -- 
    rr_4649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(117), ack => type_cast_727_inst_req_0); -- 
    -- CP-element group 118:  transition  input  no-bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Sample/ra
      -- 
    ra_4650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => send_output_CP_3660_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  no-bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	115 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_727_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Sample/rr
      -- 
    ca_4655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => send_output_CP_3660_elements(119)); -- 
    rr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(119), ack => type_cast_728_inst_req_0); -- 
    -- CP-element group 120:  transition  input  no-bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Sample/ra
      -- 
    ra_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_0, ack => send_output_CP_3660_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  no-bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	115 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (27) 
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/type_cast_728_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_offset_calculated
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_resized_0
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_scaled_0
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_computed_0
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_resize_0/$entry
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_resize_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_resize_0/index_resize_req
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_resize_0/index_resize_ack
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_scale_0/$entry
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_scale_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_scale_0/scale_rename_req
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_index_scale_0/scale_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_final_index_sum_regn/$entry
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_final_index_sum_regn/$exit
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_final_index_sum_regn/req
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_final_index_sum_regn/ack
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/array_obj_ref_732_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_request/$entry
      -- CP-element group 121: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_request/req
      -- 
    ca_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_1, ack => send_output_CP_3660_elements(121)); -- 
    req_4698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(121), ack => addr_of_733_final_reg_req_0); -- 
    -- CP-element group 122:  transition  input  no-bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	133 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_request/$exit
      -- CP-element group 122: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_request/ack
      -- 
    ack_4699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_733_final_reg_ack_0, ack => send_output_CP_3660_elements(122)); -- 
    -- CP-element group 123:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	115 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (24) 
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_complete/$exit
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/addr_of_733_complete/ack
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_word_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_root_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_address_resized
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_addr_resize/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_addr_resize/$exit
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_addr_resize/base_resize_req
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_addr_resize/base_resize_ack
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_plus_offset/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_plus_offset/$exit
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_plus_offset/sum_rename_req
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_base_plus_offset/sum_rename_ack
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_word_addrgen/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_word_addrgen/$exit
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_word_addrgen/root_register_req
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_word_addrgen/root_register_ack
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/word_0/rr
      -- 
    ack_4704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_733_final_reg_ack_1, ack => send_output_CP_3660_elements(123)); -- 
    rr_4737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(123), ack => ptr_deref_737_load_0_req_0); -- 
    -- CP-element group 124:  transition  input  no-bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Sample/word_access_start/word_0/ra
      -- 
    ra_4738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_737_load_0_ack_0, ack => send_output_CP_3660_elements(124)); -- 
    -- CP-element group 125:  transition  input  no-bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	115 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/word_access_complete/word_0/ca
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/ptr_deref_737_Merge/$entry
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/ptr_deref_737_Merge/$exit
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/ptr_deref_737_Merge/merge_req
      -- CP-element group 125: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_737_Update/ptr_deref_737_Merge/merge_ack
      -- 
    ca_4749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_737_load_0_ack_1, ack => send_output_CP_3660_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  no-bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	115 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (9) 
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/ptr_deref_740_Split/$entry
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/ptr_deref_740_Split/$exit
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/ptr_deref_740_Split/split_req
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/ptr_deref_740_Split/split_ack
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/$entry
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/word_0/rr
      -- 
    rr_4792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(126), ack => ptr_deref_740_store_0_req_0); -- 
    send_output_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(115) & send_output_CP_3660_elements(125);
      gj_send_output_cp_element_group_126 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  no-bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	132 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/$exit
      -- CP-element group 127: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/word_0/$exit
      -- CP-element group 127: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Sample/word_access_start/word_0/ra
      -- 
    ra_4793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_740_store_0_ack_0, ack => send_output_CP_3660_elements(127)); -- 
    -- CP-element group 128:  transition  input  no-bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	115 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	133 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_Update/word_access_complete/word_0/ca
      -- 
    ca_4804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_740_store_0_ack_1, ack => send_output_CP_3660_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  no-bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	115 
    -- CP-element group 129: 	132 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/$entry
      -- CP-element group 129: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/word_0/$entry
      -- CP-element group 129: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/word_0/rr
      -- 
    rr_4837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(129), ack => ptr_deref_745_load_0_req_0); -- 
    send_output_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(115) & send_output_CP_3660_elements(132);
      gj_send_output_cp_element_group_129 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  no-bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/$exit
      -- CP-element group 130: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/word_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Sample/word_access_start/word_0/ra
      -- 
    ra_4838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_745_load_0_ack_0, ack => send_output_CP_3660_elements(130)); -- 
    -- CP-element group 131:  transition  input  no-bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	115 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/$exit
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/word_0/$exit
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/word_access_complete/word_0/ca
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/ptr_deref_745_Merge/$entry
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/ptr_deref_745_Merge/$exit
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/ptr_deref_745_Merge/merge_req
      -- CP-element group 131: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_745_Update/ptr_deref_745_Merge/merge_ack
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_745_load_0_ack_1, ack => send_output_CP_3660_elements(131)); -- 
    -- CP-element group 132:  transition  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	127 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	129 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/ptr_deref_740_ptr_deref_745_delay
      -- 
    -- Element group send_output_CP_3660_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(127), ack => send_output_CP_3660_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	122 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	15 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_566/assign_stmt_724_to_assign_stmt_746/$exit
      -- 
    send_output_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(122) & send_output_CP_3660_elements(128) & send_output_CP_3660_elements(131);
      gj_send_output_cp_element_group_133 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	15 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_566/assign_stmt_749/$entry
      -- CP-element group 134: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Sample/req
      -- 
    req_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(134), ack => WPIPE_code_block_out_747_inst_req_0); -- 
    send_output_CP_3660_elements(134) <= send_output_CP_3660_elements(15);
    -- CP-element group 135:  transition  input  output  no-bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_update_start_
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Sample/ack
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Update/req
      -- 
    ack_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_code_block_out_747_inst_ack_0, ack => send_output_CP_3660_elements(135)); -- 
    req_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(135), ack => WPIPE_code_block_out_747_inst_req_1); -- 
    -- CP-element group 136:  transition  input  no-bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	16 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_566/assign_stmt_749/$exit
      -- CP-element group 136: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_566/assign_stmt_749/WPIPE_code_block_out_747_Update/ack
      -- 
    ack_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_code_block_out_747_inst_ack_1, ack => send_output_CP_3660_elements(136)); -- 
    -- CP-element group 137:  join  fork  transition  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	17 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	141 
    -- CP-element group 137: 	142 
    -- CP-element group 137: 	144 
    -- CP-element group 137:  members (51) 
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_update_start_
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_word_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_root_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_address_resized
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_addr_resize/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_addr_resize/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_addr_resize/base_resize_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_addr_resize/base_resize_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_plus_offset/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_plus_offset/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_plus_offset/sum_rename_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_base_plus_offset/sum_rename_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_word_addrgen/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_word_addrgen/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_word_addrgen/root_register_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_word_addrgen/root_register_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/word_0/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/word_0/rr
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/word_0/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/word_0/cr
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_update_start_
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_update_start_
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_word_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_root_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_address_resized
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_addr_resize/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_addr_resize/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_addr_resize/base_resize_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_addr_resize/base_resize_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_plus_offset/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_plus_offset/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_plus_offset/sum_rename_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_base_plus_offset/sum_rename_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_word_addrgen/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_word_addrgen/$exit
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_word_addrgen/root_register_req
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_word_addrgen/root_register_ack
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/word_0/$entry
      -- CP-element group 137: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/word_0/cr
      -- 
    cr_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(137), ack => ptr_deref_754_load_0_req_1); -- 
    rr_4908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(137), ack => ptr_deref_754_load_0_req_0); -- 
    cr_4938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(137), ack => ADD_u32_u32_760_inst_req_1); -- 
    cr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(137), ack => ptr_deref_763_store_0_req_1); -- 
    send_output_CP_3660_elements(137) <= send_output_CP_3660_elements(17);
    -- CP-element group 138:  transition  input  no-bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	145 
    -- CP-element group 138:  members (5) 
      -- CP-element group 138: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/$exit
      -- CP-element group 138: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/word_0/$exit
      -- CP-element group 138: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Sample/word_access_start/word_0/ra
      -- 
    ra_4909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_754_load_0_ack_0, ack => send_output_CP_3660_elements(138)); -- 
    -- CP-element group 139:  transition  input  output  no-bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/$exit
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/word_0/$exit
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/word_access_complete/word_0/ca
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/ptr_deref_754_Merge/$entry
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/ptr_deref_754_Merge/$exit
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/ptr_deref_754_Merge/merge_req
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_Update/ptr_deref_754_Merge/merge_ack
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Sample/rr
      -- 
    ca_4920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_754_load_0_ack_1, ack => send_output_CP_3660_elements(139)); -- 
    rr_4933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(139), ack => ADD_u32_u32_760_inst_req_0); -- 
    -- CP-element group 140:  transition  input  no-bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Sample/ra
      -- 
    ra_4934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_760_inst_ack_0, ack => send_output_CP_3660_elements(140)); -- 
    -- CP-element group 141:  transition  input  no-bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	137 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ADD_u32_u32_760_Update/ca
      -- 
    ca_4939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_760_inst_ack_1, ack => send_output_CP_3660_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  no-bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	137 
    -- CP-element group 142: 	141 
    -- CP-element group 142: 	145 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/ptr_deref_763_Split/$entry
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/ptr_deref_763_Split/$exit
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/ptr_deref_763_Split/split_req
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/ptr_deref_763_Split/split_ack
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/word_0/rr
      -- 
    rr_4977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(142), ack => ptr_deref_763_store_0_req_0); -- 
    send_output_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(137) & send_output_CP_3660_elements(141) & send_output_CP_3660_elements(145);
      gj_send_output_cp_element_group_142 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  no-bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/$exit
      -- CP-element group 143: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Sample/word_access_start/word_0/ra
      -- 
    ra_4978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_763_store_0_ack_0, ack => send_output_CP_3660_elements(143)); -- 
    -- CP-element group 144:  transition  input  no-bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	137 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	18 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/$exit
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/$exit
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_763_Update/word_access_complete/word_0/ca
      -- 
    ca_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_763_store_0_ack_1, ack => send_output_CP_3660_elements(144)); -- 
    -- CP-element group 145:  transition  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	138 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	142 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_566/assign_stmt_755_to_assign_stmt_765/ptr_deref_754_ptr_deref_763_delay
      -- 
    -- Element group send_output_CP_3660_elements(145) is a control-delay.
    cp_element_145_delay: control_delay_element  generic map(name => " 145_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(138), ack => send_output_CP_3660_elements(145), clk => clk, reset =>reset);
    -- CP-element group 146:  join  fork  transition  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	19 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (31) 
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_update_start_
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_address_calculated
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_word_address_calculated
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_root_address_calculated
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_address_resized
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_addr_resize/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_addr_resize/$exit
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_addr_resize/base_resize_req
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_addr_resize/base_resize_ack
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_plus_offset/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_plus_offset/$exit
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_plus_offset/sum_rename_req
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_base_plus_offset/sum_rename_ack
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_word_addrgen/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_word_addrgen/$exit
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_word_addrgen/root_register_req
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_word_addrgen/root_register_ack
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/ptr_deref_769_Split/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/ptr_deref_769_Split/$exit
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/ptr_deref_769_Split/split_req
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/ptr_deref_769_Split/split_ack
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/word_0/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/word_0/rr
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/word_0/$entry
      -- CP-element group 146: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/word_0/cr
      -- 
    cr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(146), ack => ptr_deref_769_store_0_req_1); -- 
    rr_5031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(146), ack => ptr_deref_769_store_0_req_0); -- 
    send_output_CP_3660_elements(146) <= send_output_CP_3660_elements(19);
    -- CP-element group 147:  transition  input  no-bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/$exit
      -- CP-element group 147: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/word_0/$exit
      -- CP-element group 147: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Sample/word_access_start/word_0/ra
      -- 
    ra_5032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_769_store_0_ack_0, ack => send_output_CP_3660_elements(147)); -- 
    -- CP-element group 148:  transition  input  no-bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	20 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/$exit
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/$exit
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/word_0/$exit
      -- CP-element group 148: 	 branch_block_stmt_566/assign_stmt_772/ptr_deref_769_Update/word_access_complete/word_0/ca
      -- 
    ca_5043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_769_store_0_ack_1, ack => send_output_CP_3660_elements(148)); -- 
    -- CP-element group 149:  join  fork  transition  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	21 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	152 
    -- CP-element group 149: 	153 
    -- CP-element group 149: 	155 
    -- CP-element group 149: 	158 
    -- CP-element group 149:  members (45) 
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_update_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_word_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_root_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_address_resized
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_addr_resize/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_addr_resize/$exit
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_addr_resize/base_resize_req
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_addr_resize/base_resize_ack
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_plus_offset/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_plus_offset/$exit
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_plus_offset/sum_rename_req
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_base_plus_offset/sum_rename_ack
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_word_addrgen/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_word_addrgen/$exit
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_word_addrgen/root_register_req
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_word_addrgen/root_register_ack
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/word_0/rr
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/word_0/cr
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_update_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_word_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_root_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/word_0/rr
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/word_0/cr
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_update_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_update_start_
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Update/cr
      -- 
    cr_5090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => ptr_deref_777_load_0_req_1); -- 
    rr_5079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => ptr_deref_777_load_0_req_0); -- 
    cr_5123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => LOAD_ncols_780_load_0_req_1); -- 
    rr_5112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => LOAD_ncols_780_load_0_req_0); -- 
    cr_5142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => type_cast_784_inst_req_1); -- 
    cr_5156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(149), ack => SLT_i32_u1_791_inst_req_1); -- 
    send_output_CP_3660_elements(149) <= send_output_CP_3660_elements(21);
    -- CP-element group 150:  transition  input  no-bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/$exit
      -- CP-element group 150: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/word_0/$exit
      -- CP-element group 150: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Sample/word_access_start/word_0/ra
      -- 
    ra_5080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_777_load_0_ack_0, ack => send_output_CP_3660_elements(150)); -- 
    -- CP-element group 151:  transition  input  no-bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/$exit
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/word_0/$exit
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/word_access_complete/word_0/ca
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/ptr_deref_777_Merge/$entry
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/ptr_deref_777_Merge/$exit
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/ptr_deref_777_Merge/merge_req
      -- CP-element group 151: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/ptr_deref_777_Update/ptr_deref_777_Merge/merge_ack
      -- 
    ca_5091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_777_load_0_ack_1, ack => send_output_CP_3660_elements(151)); -- 
    -- CP-element group 152:  transition  input  no-bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	149 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (5) 
      -- CP-element group 152: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/$exit
      -- CP-element group 152: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/word_0/$exit
      -- CP-element group 152: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Sample/word_access_start/word_0/ra
      -- 
    ra_5113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_780_load_0_ack_0, ack => send_output_CP_3660_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  no-bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	149 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (12) 
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/$exit
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/word_0/$exit
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/word_access_complete/word_0/ca
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/LOAD_ncols_780_Merge/$entry
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/LOAD_ncols_780_Merge/$exit
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/LOAD_ncols_780_Merge/merge_req
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/LOAD_ncols_780_Update/LOAD_ncols_780_Merge/merge_ack
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Sample/rr
      -- 
    ca_5124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_780_load_0_ack_1, ack => send_output_CP_3660_elements(153)); -- 
    rr_5137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(153), ack => type_cast_784_inst_req_0); -- 
    -- CP-element group 154:  transition  input  no-bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Sample/ra
      -- 
    ra_5138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_0, ack => send_output_CP_3660_elements(154)); -- 
    -- CP-element group 155:  transition  input  no-bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	149 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/type_cast_784_Update/ca
      -- 
    ca_5143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_1, ack => send_output_CP_3660_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Sample/rr
      -- 
    rr_5151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(156), ack => SLT_i32_u1_791_inst_req_0); -- 
    send_output_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(151) & send_output_CP_3660_elements(155);
      gj_send_output_cp_element_group_156 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  no-bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Sample/ra
      -- 
    ra_5152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_791_inst_ack_0, ack => send_output_CP_3660_elements(157)); -- 
    -- CP-element group 158:  transition  input  no-bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	149 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	22 
    -- CP-element group 158:  members (4) 
      -- CP-element group 158: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/$exit
      -- CP-element group 158: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_566/assign_stmt_778_to_assign_stmt_792/SLT_i32_u1_791_Update/ca
      -- 
    ca_5157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_791_inst_ack_1, ack => send_output_CP_3660_elements(158)); -- 
    -- CP-element group 159:  transition  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	22 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_566/if_stmt_793_dead_link/$entry
      -- 
    send_output_CP_3660_elements(159) <= send_output_CP_3660_elements(22);
    -- CP-element group 160:  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	22 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_566/if_stmt_793_eval_test/$entry
      -- CP-element group 160: 	 branch_block_stmt_566/if_stmt_793_eval_test/$exit
      -- CP-element group 160: 	 branch_block_stmt_566/if_stmt_793_eval_test/branch_req
      -- 
    branch_req_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(160), ack => if_stmt_793_branch_req_0); -- 
    send_output_CP_3660_elements(160) <= send_output_CP_3660_elements(22);
    -- CP-element group 161:  branch  place  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	164 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_566/R_iNsTr_52_794_place
      -- 
    send_output_CP_3660_elements(161) <= send_output_CP_3660_elements(160);
    -- CP-element group 162:  transition  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_566/if_stmt_793_if_link/$entry
      -- 
    send_output_CP_3660_elements(162) <= send_output_CP_3660_elements(161);
    -- CP-element group 163:  transition  input  no-bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_566/if_stmt_793_if_link/$exit
      -- CP-element group 163: 	 branch_block_stmt_566/if_stmt_793_if_link/if_choice_transition
      -- 
    if_choice_transition_5170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_793_branch_ack_1, ack => send_output_CP_3660_elements(163)); -- 
    -- CP-element group 164:  transition  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_566/if_stmt_793_else_link/$entry
      -- 
    send_output_CP_3660_elements(164) <= send_output_CP_3660_elements(161);
    -- CP-element group 165:  transition  input  no-bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_566/if_stmt_793_else_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_566/if_stmt_793_else_link/else_choice_transition
      -- 
    else_choice_transition_5174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_793_branch_ack_0, ack => send_output_CP_3660_elements(165)); -- 
    -- CP-element group 166:  place  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	163 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	232 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_566/bb_9_bb_10
      -- 
    send_output_CP_3660_elements(166) <= send_output_CP_3660_elements(163);
    -- CP-element group 167:  place  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	238 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_566/bb_9_bb_12
      -- 
    send_output_CP_3660_elements(167) <= send_output_CP_3660_elements(165);
    -- CP-element group 168:  join  fork  transition  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	23 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: 	170 
    -- CP-element group 168: 	172 
    -- CP-element group 168: 	174 
    -- CP-element group 168: 	176 
    -- CP-element group 168: 	178 
    -- CP-element group 168: 	179 
    -- CP-element group 168: 	181 
    -- CP-element group 168: 	182 
    -- CP-element group 168: 	184 
    -- CP-element group 168:  members (83) 
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_word_addrgen/root_register_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_word_addrgen/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/word_0/cr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_complete/req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_word_addrgen/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_word_addrgen/root_register_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_word_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_addr_resize/base_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_addr_resize/base_resize_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_addr_resize/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_addr_resize/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_base_address_resized
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_word_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_address_resized
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_addr_resize/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_addr_resize/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_addr_resize/base_resize_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_addr_resize/base_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_word_addrgen/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_word_addrgen/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_word_addrgen/root_register_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_word_addrgen/root_register_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/word_0/rr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/word_0/cr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/word_0/cr
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_update_start_
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_word_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_address_resized
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_addr_resize/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_addr_resize/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_addr_resize/base_resize_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_addr_resize/base_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_word_addrgen/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_word_addrgen/$exit
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_word_addrgen/root_register_req
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_word_addrgen/root_register_ack
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/word_0/cr
      -- 
    cr_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => ptr_deref_802_load_0_req_1); -- 
    rr_5212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => ptr_deref_802_load_0_req_0); -- 
    cr_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => type_cast_807_inst_req_1); -- 
    cr_5246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => type_cast_806_inst_req_1); -- 
    req_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => addr_of_812_final_reg_req_1); -- 
    cr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => ptr_deref_816_load_0_req_1); -- 
    cr_5395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => ptr_deref_819_store_0_req_1); -- 
    cr_5440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(168), ack => ptr_deref_824_load_0_req_1); -- 
    send_output_CP_3660_elements(168) <= send_output_CP_3660_elements(23);
    -- CP-element group 169:  transition  input  no-bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/$exit
      -- CP-element group 169: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/word_0/$exit
      -- CP-element group 169: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Sample/word_access_start/word_0/ra
      -- 
    ra_5213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_802_load_0_ack_0, ack => send_output_CP_3660_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  no-bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (12) 
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/word_0/$exit
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/word_access_complete/word_0/ca
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/ptr_deref_802_Merge/$entry
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/ptr_deref_802_Merge/$exit
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/ptr_deref_802_Merge/merge_req
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_802_Update/ptr_deref_802_Merge/merge_ack
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Sample/rr
      -- 
    ca_5224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_802_load_0_ack_1, ack => send_output_CP_3660_elements(170)); -- 
    rr_5241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(170), ack => type_cast_806_inst_req_0); -- 
    -- CP-element group 171:  transition  input  no-bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Sample/ra
      -- 
    ra_5242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_0, ack => send_output_CP_3660_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  no-bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	168 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_806_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Sample/rr
      -- 
    ca_5247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_1, ack => send_output_CP_3660_elements(172)); -- 
    rr_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(172), ack => type_cast_807_inst_req_0); -- 
    -- CP-element group 173:  transition  input  no-bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Sample/ra
      -- 
    ra_5252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => send_output_CP_3660_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  no-bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	168 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (27) 
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_request/req
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_request/$entry
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/type_cast_807_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_offset_calculated
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_resized_0
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_scaled_0
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_computed_0
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_resize_0/$entry
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_resize_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_resize_0/index_resize_req
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_resize_0/index_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_scale_0/$entry
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_scale_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_scale_0/scale_rename_req
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_index_scale_0/scale_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_final_index_sum_regn/$entry
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_final_index_sum_regn/$exit
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_final_index_sum_regn/req
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_final_index_sum_regn/ack
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/array_obj_ref_811_base_plus_offset/sum_rename_ack
      -- 
    ca_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_1, ack => send_output_CP_3660_elements(174)); -- 
    req_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(174), ack => addr_of_812_final_reg_req_0); -- 
    -- CP-element group 175:  transition  input  no-bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	186 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_request/ack
      -- CP-element group 175: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_request/$exit
      -- CP-element group 175: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_sample_completed_
      -- 
    ack_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_812_final_reg_ack_0, ack => send_output_CP_3660_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	168 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (24) 
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_word_address_calculated
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_address_resized
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_addr_resize/$exit
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_address_calculated
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_complete/$exit
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_root_address_calculated
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_addr_resize/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/word_0/rr
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/word_0/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_word_addrgen/root_register_ack
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_word_addrgen/root_register_req
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_word_addrgen/$exit
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_word_addrgen/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_complete/ack
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_plus_offset/sum_rename_ack
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_plus_offset/sum_rename_req
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_plus_offset/$exit
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_plus_offset/$entry
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_addr_resize/base_resize_ack
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_base_addr_resize/base_resize_req
      -- CP-element group 176: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/addr_of_812_update_completed_
      -- 
    ack_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_812_final_reg_ack_1, ack => send_output_CP_3660_elements(176)); -- 
    rr_5329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(176), ack => ptr_deref_816_load_0_req_0); -- 
    -- CP-element group 177:  transition  input  no-bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/word_0/ra
      -- CP-element group 177: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/word_0/$exit
      -- CP-element group 177: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/word_access_start/$exit
      -- CP-element group 177: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Sample/$exit
      -- 
    ra_5330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_load_0_ack_0, ack => send_output_CP_3660_elements(177)); -- 
    -- CP-element group 178:  transition  input  no-bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	168 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/word_0/ca
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/ptr_deref_816_Merge/$entry
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/ptr_deref_816_Merge/$exit
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/ptr_deref_816_Merge/merge_req
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/ptr_deref_816_Merge/merge_ack
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/word_0/$exit
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/word_access_complete/$exit
      -- CP-element group 178: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_816_Update/$exit
      -- 
    ca_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_load_0_ack_1, ack => send_output_CP_3660_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  no-bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	168 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/ptr_deref_819_Split/$entry
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/ptr_deref_819_Split/$exit
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/ptr_deref_819_Split/split_req
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/ptr_deref_819_Split/split_ack
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/$entry
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/word_0/$entry
      -- CP-element group 179: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/word_0/rr
      -- 
    rr_5384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(179), ack => ptr_deref_819_store_0_req_0); -- 
    send_output_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(168) & send_output_CP_3660_elements(178);
      gj_send_output_cp_element_group_179 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  transition  input  no-bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	185 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/$exit
      -- CP-element group 180: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/word_0/$exit
      -- CP-element group 180: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Sample/word_access_start/word_0/ra
      -- 
    ra_5385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_store_0_ack_0, ack => send_output_CP_3660_elements(180)); -- 
    -- CP-element group 181:  transition  input  no-bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	168 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_Update/word_access_complete/word_0/ca
      -- 
    ca_5396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_store_0_ack_1, ack => send_output_CP_3660_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  no-bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	168 
    -- CP-element group 182: 	185 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/$entry
      -- CP-element group 182: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/word_0/$entry
      -- CP-element group 182: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/word_0/rr
      -- 
    rr_5429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(182), ack => ptr_deref_824_load_0_req_0); -- 
    send_output_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(168) & send_output_CP_3660_elements(185);
      gj_send_output_cp_element_group_182 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  transition  input  no-bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/$exit
      -- CP-element group 183: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/word_0/$exit
      -- CP-element group 183: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Sample/word_access_start/word_0/ra
      -- 
    ra_5430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_824_load_0_ack_0, ack => send_output_CP_3660_elements(183)); -- 
    -- CP-element group 184:  transition  input  no-bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	168 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/$exit
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/word_0/$exit
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/word_access_complete/word_0/ca
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/ptr_deref_824_Merge/$entry
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/ptr_deref_824_Merge/$exit
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/ptr_deref_824_Merge/merge_req
      -- CP-element group 184: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_824_Update/ptr_deref_824_Merge/merge_ack
      -- 
    ca_5441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_824_load_0_ack_1, ack => send_output_CP_3660_elements(184)); -- 
    -- CP-element group 185:  transition  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	180 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	182 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/ptr_deref_819_ptr_deref_824_delay
      -- 
    -- Element group send_output_CP_3660_elements(185) is a control-delay.
    cp_element_185_delay: control_delay_element  generic map(name => " 185_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(180), ack => send_output_CP_3660_elements(185), clk => clk, reset =>reset);
    -- CP-element group 186:  join  transition  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	175 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	24 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_566/assign_stmt_803_to_assign_stmt_825/$exit
      -- 
    send_output_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(175) & send_output_CP_3660_elements(181) & send_output_CP_3660_elements(184);
      gj_send_output_cp_element_group_186 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  transition  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	24 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (4) 
      -- CP-element group 187: 	 branch_block_stmt_566/assign_stmt_828/$entry
      -- CP-element group 187: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Sample/req
      -- 
    req_5458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(187), ack => WPIPE_aPriori_out_826_inst_req_0); -- 
    send_output_CP_3660_elements(187) <= send_output_CP_3660_elements(24);
    -- CP-element group 188:  transition  input  output  no-bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (6) 
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_update_start_
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Sample/ack
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Update/req
      -- 
    ack_5459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_aPriori_out_826_inst_ack_0, ack => send_output_CP_3660_elements(188)); -- 
    req_5463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(188), ack => WPIPE_aPriori_out_826_inst_req_1); -- 
    -- CP-element group 189:  transition  input  no-bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	25 
    -- CP-element group 189:  members (4) 
      -- CP-element group 189: 	 branch_block_stmt_566/assign_stmt_828/$exit
      -- CP-element group 189: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_566/assign_stmt_828/WPIPE_aPriori_out_826_Update/ack
      -- 
    ack_5464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_aPriori_out_826_inst_ack_1, ack => send_output_CP_3660_elements(189)); -- 
    -- CP-element group 190:  join  fork  transition  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	26 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	194 
    -- CP-element group 190: 	195 
    -- CP-element group 190: 	197 
    -- CP-element group 190:  members (51) 
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_update_start_
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_word_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_root_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_address_resized
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_addr_resize/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_addr_resize/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_addr_resize/base_resize_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_addr_resize/base_resize_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_plus_offset/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_plus_offset/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_plus_offset/sum_rename_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_base_plus_offset/sum_rename_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_word_addrgen/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_word_addrgen/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_word_addrgen/root_register_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_word_addrgen/root_register_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/word_0/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/word_0/rr
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/word_0/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/word_0/cr
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_update_start_
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_update_start_
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_word_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_root_address_calculated
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_address_resized
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_addr_resize/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_addr_resize/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_addr_resize/base_resize_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_addr_resize/base_resize_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_plus_offset/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_plus_offset/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_plus_offset/sum_rename_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_base_plus_offset/sum_rename_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_word_addrgen/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_word_addrgen/$exit
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_word_addrgen/root_register_req
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_word_addrgen/root_register_ack
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/word_0/$entry
      -- CP-element group 190: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/word_0/cr
      -- 
    cr_5511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(190), ack => ptr_deref_833_load_0_req_1); -- 
    rr_5500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(190), ack => ptr_deref_833_load_0_req_0); -- 
    cr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(190), ack => ADD_u32_u32_839_inst_req_1); -- 
    cr_5580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(190), ack => ptr_deref_842_store_0_req_1); -- 
    send_output_CP_3660_elements(190) <= send_output_CP_3660_elements(26);
    -- CP-element group 191:  transition  input  no-bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	198 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/$exit
      -- CP-element group 191: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/word_0/$exit
      -- CP-element group 191: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Sample/word_access_start/word_0/ra
      -- 
    ra_5501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_load_0_ack_0, ack => send_output_CP_3660_elements(191)); -- 
    -- CP-element group 192:  transition  input  output  no-bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (12) 
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/$exit
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/word_0/$exit
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/word_access_complete/word_0/ca
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/ptr_deref_833_Merge/$entry
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/ptr_deref_833_Merge/$exit
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/ptr_deref_833_Merge/merge_req
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_Update/ptr_deref_833_Merge/merge_ack
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Sample/rr
      -- 
    ca_5512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_load_0_ack_1, ack => send_output_CP_3660_elements(192)); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(192), ack => ADD_u32_u32_839_inst_req_0); -- 
    -- CP-element group 193:  transition  input  no-bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Sample/ra
      -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_839_inst_ack_0, ack => send_output_CP_3660_elements(193)); -- 
    -- CP-element group 194:  transition  input  no-bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ADD_u32_u32_839_Update/ca
      -- 
    ca_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_839_inst_ack_1, ack => send_output_CP_3660_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  no-bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	190 
    -- CP-element group 195: 	194 
    -- CP-element group 195: 	198 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/ptr_deref_842_Split/$entry
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/ptr_deref_842_Split/$exit
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/ptr_deref_842_Split/split_req
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/ptr_deref_842_Split/split_ack
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/$entry
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/word_0/$entry
      -- CP-element group 195: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/word_0/rr
      -- 
    rr_5569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(195), ack => ptr_deref_842_store_0_req_0); -- 
    send_output_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 32) := "send_output_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= send_output_CP_3660_elements(190) & send_output_CP_3660_elements(194) & send_output_CP_3660_elements(198);
      gj_send_output_cp_element_group_195 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => send_output_CP_3660_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  transition  input  no-bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/$exit
      -- CP-element group 196: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/word_0/$exit
      -- CP-element group 196: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Sample/word_access_start/word_0/ra
      -- 
    ra_5570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_842_store_0_ack_0, ack => send_output_CP_3660_elements(196)); -- 
    -- CP-element group 197:  transition  input  no-bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	190 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	27 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/$exit
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/$exit
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_842_Update/word_access_complete/word_0/ca
      -- 
    ca_5581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_842_store_0_ack_1, ack => send_output_CP_3660_elements(197)); -- 
    -- CP-element group 198:  transition  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	191 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	195 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_566/assign_stmt_834_to_assign_stmt_844/ptr_deref_833_ptr_deref_842_delay
      -- 
    -- Element group send_output_CP_3660_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => send_output_CP_3660_elements(191), ack => send_output_CP_3660_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  join  fork  transition  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	28 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (27) 
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_update_start_
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_word_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_root_address_calculated
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_address_resized
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_addr_resize/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_addr_resize/$exit
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_addr_resize/base_resize_req
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_addr_resize/base_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_plus_offset/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_plus_offset/$exit
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_plus_offset/sum_rename_req
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_base_plus_offset/sum_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_word_addrgen/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_word_addrgen/$exit
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_word_addrgen/root_register_req
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_word_addrgen/root_register_ack
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/word_0/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/word_0/rr
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/word_0/$entry
      -- CP-element group 199: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/word_0/cr
      -- 
    cr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(199), ack => ptr_deref_849_load_0_req_1); -- 
    rr_5618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => send_output_CP_3660_elements(199), ack => ptr_deref_849_load_0_req_0); -- 
    send_output_CP_3660_elements(199) <= send_output_CP_3660_elements(28);
    -- CP-element group 200:  transition  input  no-bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (5) 
      -- CP-element group 200: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/$exit
      -- CP-element group 200: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/word_0/$exit
      -- CP-element group 200: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Sample/word_access_start/word_0/ra
      -- 
    ra_5619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_849_load_0_ack_0, ack => send_output_CP_3660_elements(200)); -- 
    -- CP-element group 201:  transition  input  no-bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	29 
    -- CP-element group 201:  members (10) 
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/$exit
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/$exit
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/word_0/$exit
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/word_access_complete/word_0/ca
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/ptr_deref_849_Merge/$entry
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/ptr_deref_849_Merge/$exit
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/ptr_deref_849_Merge/merge_req
      -- CP-element group 201: 	 branch_block_stmt_566/assign_stmt_850/ptr_deref_849_Update/ptr_deref_849_Merge/merge_ack
      -- 
    ca_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_849_load_0_ack_1, ack => send_output_CP_3660_elements(201)); -- 
    -- CP-element group 202:  transition  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	2 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_566/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 202: 	 branch_block_stmt_566/bb_0_bb_1_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(202) <= send_output_CP_3660_elements(2);
    -- CP-element group 203:  transition  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_566/bb_3_bb_1_PhiReq/$entry
      -- CP-element group 203: 	 branch_block_stmt_566/bb_3_bb_1_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(203) <= send_output_CP_3660_elements(9);
    -- CP-element group 204:  merge  place  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_566/merge_stmt_598_PhiReqMerge
      -- 
    send_output_CP_3660_elements(204) <= OrReduce(send_output_CP_3660_elements(202) & send_output_CP_3660_elements(203));
    -- CP-element group 205:  transition  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	3 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_566/merge_stmt_598_PhiAck/$entry
      -- CP-element group 205: 	 branch_block_stmt_566/merge_stmt_598_PhiAck/$exit
      -- CP-element group 205: 	 branch_block_stmt_566/merge_stmt_598_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(205) <= send_output_CP_3660_elements(204);
    -- CP-element group 206:  transition  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	60 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_566/bb_1_bb_2_PhiReq/$entry
      -- CP-element group 206: 	 branch_block_stmt_566/bb_1_bb_2_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(206) <= send_output_CP_3660_elements(60);
    -- CP-element group 207:  place  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_566/merge_stmt_641_PhiReqMerge
      -- 
    send_output_CP_3660_elements(207) <= send_output_CP_3660_elements(206);
    -- CP-element group 208:  transition  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	5 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_566/merge_stmt_641_PhiAck/$entry
      -- CP-element group 208: 	 branch_block_stmt_566/merge_stmt_641_PhiAck/$exit
      -- CP-element group 208: 	 branch_block_stmt_566/merge_stmt_641_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(208) <= send_output_CP_3660_elements(207);
    -- CP-element group 209:  transition  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	7 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_566/bb_2_bb_3_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_566/bb_2_bb_3_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(209) <= send_output_CP_3660_elements(7);
    -- CP-element group 210:  place  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_566/merge_stmt_672_PhiReqMerge
      -- 
    send_output_CP_3660_elements(210) <= send_output_CP_3660_elements(209);
    -- CP-element group 211:  transition  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	8 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_566/merge_stmt_672_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_566/merge_stmt_672_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_566/merge_stmt_672_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(211) <= send_output_CP_3660_elements(210);
    -- CP-element group 212:  transition  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	61 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_566/bb_1_bb_4_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_566/bb_1_bb_4_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(212) <= send_output_CP_3660_elements(61);
    -- CP-element group 213:  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_566/merge_stmt_688_PhiReqMerge
      -- 
    send_output_CP_3660_elements(213) <= send_output_CP_3660_elements(212);
    -- CP-element group 214:  transition  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	10 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_566/merge_stmt_688_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_566/merge_stmt_688_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_566/merge_stmt_688_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(214) <= send_output_CP_3660_elements(213);
    -- CP-element group 215:  transition  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	11 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_566/bb_4_bb_5_PhiReq/$entry
      -- CP-element group 215: 	 branch_block_stmt_566/bb_4_bb_5_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(215) <= send_output_CP_3660_elements(11);
    -- CP-element group 216:  transition  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	18 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_566/bb_7_bb_5_PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_566/bb_7_bb_5_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(216) <= send_output_CP_3660_elements(18);
    -- CP-element group 217:  merge  place  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_566/merge_stmt_695_PhiReqMerge
      -- 
    send_output_CP_3660_elements(217) <= OrReduce(send_output_CP_3660_elements(215) & send_output_CP_3660_elements(216));
    -- CP-element group 218:  transition  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	12 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_566/merge_stmt_695_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_566/merge_stmt_695_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_566/merge_stmt_695_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(218) <= send_output_CP_3660_elements(217);
    -- CP-element group 219:  transition  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	113 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (2) 
      -- CP-element group 219: 	 branch_block_stmt_566/bb_5_bb_6_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_566/bb_5_bb_6_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(219) <= send_output_CP_3660_elements(113);
    -- CP-element group 220:  place  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_566/merge_stmt_720_PhiReqMerge
      -- 
    send_output_CP_3660_elements(220) <= send_output_CP_3660_elements(219);
    -- CP-element group 221:  transition  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	14 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_566/merge_stmt_720_PhiAck/$entry
      -- CP-element group 221: 	 branch_block_stmt_566/merge_stmt_720_PhiAck/$exit
      -- CP-element group 221: 	 branch_block_stmt_566/merge_stmt_720_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(221) <= send_output_CP_3660_elements(220);
    -- CP-element group 222:  transition  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	16 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_566/bb_6_bb_7_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_566/bb_6_bb_7_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(222) <= send_output_CP_3660_elements(16);
    -- CP-element group 223:  place  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_566/merge_stmt_751_PhiReqMerge
      -- 
    send_output_CP_3660_elements(223) <= send_output_CP_3660_elements(222);
    -- CP-element group 224:  transition  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	17 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_566/merge_stmt_751_PhiAck/$entry
      -- CP-element group 224: 	 branch_block_stmt_566/merge_stmt_751_PhiAck/$exit
      -- CP-element group 224: 	 branch_block_stmt_566/merge_stmt_751_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(224) <= send_output_CP_3660_elements(223);
    -- CP-element group 225:  transition  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	114 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_566/bb_5_bb_8_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_566/bb_5_bb_8_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(225) <= send_output_CP_3660_elements(114);
    -- CP-element group 226:  place  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_566/merge_stmt_767_PhiReqMerge
      -- 
    send_output_CP_3660_elements(226) <= send_output_CP_3660_elements(225);
    -- CP-element group 227:  transition  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	19 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_566/merge_stmt_767_PhiAck/$entry
      -- CP-element group 227: 	 branch_block_stmt_566/merge_stmt_767_PhiAck/$exit
      -- CP-element group 227: 	 branch_block_stmt_566/merge_stmt_767_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(227) <= send_output_CP_3660_elements(226);
    -- CP-element group 228:  transition  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	27 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_566/bb_11_bb_9_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_566/bb_11_bb_9_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(228) <= send_output_CP_3660_elements(27);
    -- CP-element group 229:  transition  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	20 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_566/bb_8_bb_9_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_566/bb_8_bb_9_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(229) <= send_output_CP_3660_elements(20);
    -- CP-element group 230:  merge  place  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_566/merge_stmt_774_PhiReqMerge
      -- 
    send_output_CP_3660_elements(230) <= OrReduce(send_output_CP_3660_elements(228) & send_output_CP_3660_elements(229));
    -- CP-element group 231:  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	21 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_566/merge_stmt_774_PhiAck/$entry
      -- CP-element group 231: 	 branch_block_stmt_566/merge_stmt_774_PhiAck/$exit
      -- CP-element group 231: 	 branch_block_stmt_566/merge_stmt_774_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(231) <= send_output_CP_3660_elements(230);
    -- CP-element group 232:  transition  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	166 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (2) 
      -- CP-element group 232: 	 branch_block_stmt_566/bb_9_bb_10_PhiReq/$entry
      -- CP-element group 232: 	 branch_block_stmt_566/bb_9_bb_10_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(232) <= send_output_CP_3660_elements(166);
    -- CP-element group 233:  place  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_566/merge_stmt_799_PhiReqMerge
      -- 
    send_output_CP_3660_elements(233) <= send_output_CP_3660_elements(232);
    -- CP-element group 234:  transition  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	23 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_566/merge_stmt_799_PhiAck/$entry
      -- CP-element group 234: 	 branch_block_stmt_566/merge_stmt_799_PhiAck/$exit
      -- CP-element group 234: 	 branch_block_stmt_566/merge_stmt_799_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(234) <= send_output_CP_3660_elements(233);
    -- CP-element group 235:  transition  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	25 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_566/bb_10_bb_11_PhiReq/$entry
      -- CP-element group 235: 	 branch_block_stmt_566/bb_10_bb_11_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(235) <= send_output_CP_3660_elements(25);
    -- CP-element group 236:  place  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_566/merge_stmt_830_PhiReqMerge
      -- 
    send_output_CP_3660_elements(236) <= send_output_CP_3660_elements(235);
    -- CP-element group 237:  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	26 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_566/merge_stmt_830_PhiAck/$entry
      -- CP-element group 237: 	 branch_block_stmt_566/merge_stmt_830_PhiAck/$exit
      -- CP-element group 237: 	 branch_block_stmt_566/merge_stmt_830_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(237) <= send_output_CP_3660_elements(236);
    -- CP-element group 238:  transition  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	167 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_566/bb_9_bb_12_PhiReq/$entry
      -- CP-element group 238: 	 branch_block_stmt_566/bb_9_bb_12_PhiReq/$exit
      -- 
    send_output_CP_3660_elements(238) <= send_output_CP_3660_elements(167);
    -- CP-element group 239:  place  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (1) 
      -- CP-element group 239: 	 branch_block_stmt_566/merge_stmt_846_PhiReqMerge
      -- 
    send_output_CP_3660_elements(239) <= send_output_CP_3660_elements(238);
    -- CP-element group 240:  transition  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	28 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_566/merge_stmt_846_PhiAck/$entry
      -- CP-element group 240: 	 branch_block_stmt_566/merge_stmt_846_PhiAck/$exit
      -- CP-element group 240: 	 branch_block_stmt_566/merge_stmt_846_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(240) <= send_output_CP_3660_elements(239);
    -- CP-element group 241:  transition  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	29 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (2) 
      -- CP-element group 241: 	 branch_block_stmt_566/return___PhiReq/$entry
      -- CP-element group 241: 	 branch_block_stmt_566/return___PhiReq/$exit
      -- 
    send_output_CP_3660_elements(241) <= send_output_CP_3660_elements(29);
    -- CP-element group 242:  place  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_566/merge_stmt_852_PhiReqMerge
      -- 
    send_output_CP_3660_elements(242) <= send_output_CP_3660_elements(241);
    -- CP-element group 243:  transition  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	30 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_566/merge_stmt_852_PhiAck/$entry
      -- CP-element group 243: 	 branch_block_stmt_566/merge_stmt_852_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_566/merge_stmt_852_PhiAck/dummy
      -- 
    send_output_CP_3660_elements(243) <= send_output_CP_3660_elements(242);
    -- CP-element group 244:  transition  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	30 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_566/$exit
      -- CP-element group 244: 	 $exit
      -- 
    send_output_CP_3660_elements(244) <= send_output_CP_3660_elements(30);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal J_579 : std_logic_vector(31 downto 0);
    signal LOAD_ncol_ind_611_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncol_ind_611_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_701_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_701_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_780_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_780_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_nrows_604_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_nrows_604_word_address_0 : std_logic_vector(0 downto 0);
    signal R_iNsTr_14_652_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_14_652_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_35_731_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_35_731_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_56_810_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_56_810_scaled : std_logic_vector(9 downto 0);
    signal array_obj_ref_653_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_653_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_653_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_653_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_732_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_732_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_732_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_732_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_811_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_811_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_811_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_811_root_address : std_logic_vector(9 downto 0);
    signal iNsTr_0_575 : std_logic_vector(31 downto 0);
    signal iNsTr_10_634 : std_logic_vector(0 downto 0);
    signal iNsTr_13_645 : std_logic_vector(31 downto 0);
    signal iNsTr_14_650 : std_logic_vector(63 downto 0);
    signal iNsTr_15_655 : std_logic_vector(31 downto 0);
    signal iNsTr_16_659 : std_logic_vector(15 downto 0);
    signal iNsTr_18_667 : std_logic_vector(15 downto 0);
    signal iNsTr_24_676 : std_logic_vector(31 downto 0);
    signal iNsTr_25_682 : std_logic_vector(31 downto 0);
    signal iNsTr_28_699 : std_logic_vector(31 downto 0);
    signal iNsTr_29_702 : std_logic_vector(15 downto 0);
    signal iNsTr_30_706 : std_logic_vector(31 downto 0);
    signal iNsTr_31_713 : std_logic_vector(0 downto 0);
    signal iNsTr_34_724 : std_logic_vector(31 downto 0);
    signal iNsTr_35_729 : std_logic_vector(63 downto 0);
    signal iNsTr_36_734 : std_logic_vector(31 downto 0);
    signal iNsTr_37_738 : std_logic_vector(31 downto 0);
    signal iNsTr_39_746 : std_logic_vector(31 downto 0);
    signal iNsTr_3_602 : std_logic_vector(31 downto 0);
    signal iNsTr_45_755 : std_logic_vector(31 downto 0);
    signal iNsTr_46_761 : std_logic_vector(31 downto 0);
    signal iNsTr_49_778 : std_logic_vector(31 downto 0);
    signal iNsTr_4_605 : std_logic_vector(15 downto 0);
    signal iNsTr_50_781 : std_logic_vector(15 downto 0);
    signal iNsTr_51_785 : std_logic_vector(31 downto 0);
    signal iNsTr_52_792 : std_logic_vector(0 downto 0);
    signal iNsTr_55_803 : std_logic_vector(31 downto 0);
    signal iNsTr_56_808 : std_logic_vector(63 downto 0);
    signal iNsTr_57_813 : std_logic_vector(31 downto 0);
    signal iNsTr_58_817 : std_logic_vector(31 downto 0);
    signal iNsTr_5_609 : std_logic_vector(31 downto 0);
    signal iNsTr_60_825 : std_logic_vector(31 downto 0);
    signal iNsTr_66_834 : std_logic_vector(31 downto 0);
    signal iNsTr_67_840 : std_logic_vector(31 downto 0);
    signal iNsTr_6_612 : std_logic_vector(15 downto 0);
    signal iNsTr_7_616 : std_logic_vector(31 downto 0);
    signal iNsTr_8_621 : std_logic_vector(31 downto 0);
    signal iNsTr_9_627 : std_logic_vector(31 downto 0);
    signal ptr_deref_593_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_593_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_593_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_593_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_593_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_593_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_601_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_601_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_601_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_601_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_601_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_644_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_644_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_644_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_644_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_644_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_658_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_658_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_658_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_658_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_658_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_661_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_661_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_661_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_661_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_661_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_661_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_666_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_666_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_666_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_666_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_666_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_675_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_675_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_675_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_675_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_675_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_684_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_684_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_684_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_684_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_684_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_684_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_690_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_690_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_690_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_690_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_690_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_690_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_698_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_698_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_698_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_698_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_698_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_723_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_723_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_723_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_723_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_723_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_737_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_737_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_737_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_737_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_737_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_740_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_740_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_740_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_740_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_740_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_740_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_745_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_745_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_745_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_745_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_745_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_754_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_754_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_754_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_754_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_754_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_763_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_763_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_763_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_763_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_763_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_763_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_769_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_769_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_769_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_769_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_769_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_769_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_777_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_777_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_777_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_777_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_777_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_802_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_802_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_802_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_802_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_802_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_816_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_816_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_816_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_816_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_816_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_819_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_819_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_819_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_819_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_819_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_819_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_824_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_824_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_824_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_824_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_824_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_833_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_833_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_833_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_833_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_833_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_842_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_842_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_842_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_842_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_842_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_842_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_849_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_849_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_849_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_849_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_849_word_offset_0 : std_logic_vector(0 downto 0);
    signal type_cast_595_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_630_wire : std_logic_vector(31 downto 0);
    signal type_cast_632_wire : std_logic_vector(31 downto 0);
    signal type_cast_648_wire : std_logic_vector(63 downto 0);
    signal type_cast_680_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_692_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_709_wire : std_logic_vector(31 downto 0);
    signal type_cast_711_wire : std_logic_vector(31 downto 0);
    signal type_cast_727_wire : std_logic_vector(63 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_771_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_788_wire : std_logic_vector(31 downto 0);
    signal type_cast_790_wire : std_logic_vector(31 downto 0);
    signal type_cast_806_wire : std_logic_vector(63 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(31 downto 0);
    signal val1_587 : std_logic_vector(31 downto 0);
    signal val2_591 : std_logic_vector(31 downto 0);
    signal val_583 : std_logic_vector(31 downto 0);
    signal xxsend_outputxxbodyxxJ_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxsend_outputxxbodyxxiNsTr_0_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxsend_outputxxbodyxxval1_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxsend_outputxxbodyxxval2_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxsend_outputxxbodyxxval_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    J_579 <= "00000000000000000000000000000000";
    LOAD_ncol_ind_611_word_address_0 <= "0";
    LOAD_ncols_701_word_address_0 <= "0";
    LOAD_ncols_780_word_address_0 <= "0";
    LOAD_nrows_604_word_address_0 <= "0";
    array_obj_ref_653_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_653_resized_base_address <= "0000000000";
    array_obj_ref_732_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_732_resized_base_address <= "0000000000";
    array_obj_ref_811_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_811_resized_base_address <= "0000000000";
    iNsTr_0_575 <= "00000000000000000000000000000000";
    ptr_deref_593_word_offset_0 <= "0";
    ptr_deref_601_word_offset_0 <= "0";
    ptr_deref_644_word_offset_0 <= "0";
    ptr_deref_658_word_offset_0 <= "0000000000";
    ptr_deref_661_word_offset_0 <= "0";
    ptr_deref_666_word_offset_0 <= "0";
    ptr_deref_675_word_offset_0 <= "0";
    ptr_deref_684_word_offset_0 <= "0";
    ptr_deref_690_word_offset_0 <= "0";
    ptr_deref_698_word_offset_0 <= "0";
    ptr_deref_723_word_offset_0 <= "0";
    ptr_deref_737_word_offset_0 <= "0000000000";
    ptr_deref_740_word_offset_0 <= "0";
    ptr_deref_745_word_offset_0 <= "0";
    ptr_deref_754_word_offset_0 <= "0";
    ptr_deref_763_word_offset_0 <= "0";
    ptr_deref_769_word_offset_0 <= "0";
    ptr_deref_777_word_offset_0 <= "0";
    ptr_deref_802_word_offset_0 <= "0";
    ptr_deref_816_word_offset_0 <= "0000000000";
    ptr_deref_819_word_offset_0 <= "0";
    ptr_deref_824_word_offset_0 <= "0";
    ptr_deref_833_word_offset_0 <= "0";
    ptr_deref_842_word_offset_0 <= "0";
    ptr_deref_849_word_offset_0 <= "0";
    type_cast_595_wire_constant <= "00000000000000000000000000000000";
    type_cast_625_wire_constant <= "00000000000000000000000000000011";
    type_cast_680_wire_constant <= "00000000000000000000000000000001";
    type_cast_692_wire_constant <= "00000000000000000000000000000000";
    type_cast_759_wire_constant <= "00000000000000000000000000000001";
    type_cast_771_wire_constant <= "00000000000000000000000000000000";
    type_cast_838_wire_constant <= "00000000000000000000000000000001";
    val1_587 <= "00000000000000000000000000000000";
    val2_591 <= "00000000000000000000000000000000";
    val_583 <= "00000000000000000000000000000000";
    xxsend_outputxxbodyxxJ_alloc_base_address <= "0";
    xxsend_outputxxbodyxxiNsTr_0_alloc_base_address <= "0";
    xxsend_outputxxbodyxxval1_alloc_base_address <= "0";
    xxsend_outputxxbodyxxval2_alloc_base_address <= "0";
    xxsend_outputxxbodyxxval_alloc_base_address <= "0";
    addr_of_654_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_654_final_reg_req_0;
      addr_of_654_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_654_final_reg_req_1;
      addr_of_654_final_reg_ack_1<= rack(0);
      addr_of_654_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_654_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_653_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_15_655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_733_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_733_final_reg_req_0;
      addr_of_733_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_733_final_reg_req_1;
      addr_of_733_final_reg_ack_1<= rack(0);
      addr_of_733_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_733_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_732_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_36_734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_812_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_812_final_reg_req_0;
      addr_of_812_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_812_final_reg_req_1;
      addr_of_812_final_reg_ack_1<= rack(0);
      addr_of_812_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_812_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_811_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_57_813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_4_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_5_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_6_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_7_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_630_inst
    process(iNsTr_3_602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_3_602(31 downto 0);
      type_cast_630_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_632_inst
    process(iNsTr_9_627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_9_627(31 downto 0);
      type_cast_632_wire <= tmp_var; -- 
    end process;
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_648_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_705_inst_req_0;
      type_cast_705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_705_inst_req_1;
      type_cast_705_inst_ack_1<= rack(0);
      type_cast_705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_29_702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_30_706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_709_inst
    process(iNsTr_28_699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_28_699(31 downto 0);
      type_cast_709_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_711_inst
    process(iNsTr_30_706) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_30_706(31 downto 0);
      type_cast_711_wire <= tmp_var; -- 
    end process;
    type_cast_728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_728_inst_req_0;
      type_cast_728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_728_inst_req_1;
      type_cast_728_inst_ack_1<= rack(0);
      type_cast_728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_727_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_35_729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_784_inst_req_0;
      type_cast_784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_784_inst_req_1;
      type_cast_784_inst_ack_1<= rack(0);
      type_cast_784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_50_781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_51_785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_788_inst
    process(iNsTr_49_778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_49_778(31 downto 0);
      type_cast_788_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_790_inst
    process(iNsTr_51_785) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_51_785(31 downto 0);
      type_cast_790_wire <= tmp_var; -- 
    end process;
    type_cast_807_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_807_inst_req_0;
      type_cast_807_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_807_inst_req_1;
      type_cast_807_inst_ack_1<= rack(0);
      type_cast_807_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_807_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_806_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_56_808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_ncol_ind_611_gather_scatter
    process(LOAD_ncol_ind_611_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncol_ind_611_data_0;
      ov(15 downto 0) := iv;
      iNsTr_6_612 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_701_gather_scatter
    process(LOAD_ncols_701_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_701_data_0;
      ov(15 downto 0) := iv;
      iNsTr_29_702 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_780_gather_scatter
    process(LOAD_ncols_780_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_780_data_0;
      ov(15 downto 0) := iv;
      iNsTr_50_781 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_nrows_604_gather_scatter
    process(LOAD_nrows_604_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_nrows_604_data_0;
      ov(15 downto 0) := iv;
      iNsTr_4_605 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_0_rename
    process(R_iNsTr_14_652_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_14_652_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_14_652_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_0_resize
    process(iNsTr_14_650) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_14_650;
      ov := iv(9 downto 0);
      R_iNsTr_14_652_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_offset
    process(R_iNsTr_14_652_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_14_652_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_653_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_root_address_inst
    process(array_obj_ref_653_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_653_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_653_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_732_index_0_rename
    process(R_iNsTr_35_731_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_35_731_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_35_731_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_732_index_0_resize
    process(iNsTr_35_729) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_729;
      ov := iv(9 downto 0);
      R_iNsTr_35_731_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_732_index_offset
    process(R_iNsTr_35_731_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_35_731_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_732_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_732_root_address_inst
    process(array_obj_ref_732_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_732_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_732_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_index_0_rename
    process(R_iNsTr_56_810_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_56_810_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_56_810_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_index_0_resize
    process(iNsTr_56_808) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_56_808;
      ov := iv(9 downto 0);
      R_iNsTr_56_810_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_index_offset
    process(R_iNsTr_56_810_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_56_810_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_811_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_811_root_address_inst
    process(array_obj_ref_811_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_811_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_811_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_593_addr_0
    process(ptr_deref_593_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_593_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_593_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_593_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_593_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_593_gather_scatter
    process(type_cast_595_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_595_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_593_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_593_root_address_inst
    process(ptr_deref_593_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_593_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_593_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_addr_0
    process(ptr_deref_601_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_601_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_601_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_601_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_gather_scatter
    process(ptr_deref_601_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_601_data_0;
      ov(31 downto 0) := iv;
      iNsTr_3_602 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_root_address_inst
    process(ptr_deref_601_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_601_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_601_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_644_addr_0
    process(ptr_deref_644_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_644_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_644_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_644_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_644_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_644_gather_scatter
    process(ptr_deref_644_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_644_data_0;
      ov(31 downto 0) := iv;
      iNsTr_13_645 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_644_root_address_inst
    process(ptr_deref_644_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_644_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_644_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_658_addr_0
    process(ptr_deref_658_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_658_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_658_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_658_base_resize
    process(iNsTr_15_655) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_655;
      ov := iv(9 downto 0);
      ptr_deref_658_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_658_gather_scatter
    process(ptr_deref_658_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_658_data_0;
      ov(15 downto 0) := iv;
      iNsTr_16_659 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_658_root_address_inst
    process(ptr_deref_658_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_658_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_658_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_661_addr_0
    process(ptr_deref_661_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_661_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_661_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_661_base_resize
    process(val_583) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_583;
      ov := iv(0 downto 0);
      ptr_deref_661_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_661_gather_scatter
    process(iNsTr_16_659) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_659;
      ov(15 downto 0) := iv;
      ptr_deref_661_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_661_root_address_inst
    process(ptr_deref_661_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_661_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_661_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_addr_0
    process(ptr_deref_666_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_666_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_666_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_base_resize
    process(val_583) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_583;
      ov := iv(0 downto 0);
      ptr_deref_666_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_gather_scatter
    process(ptr_deref_666_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_666_data_0;
      ov(15 downto 0) := iv;
      iNsTr_18_667 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_root_address_inst
    process(ptr_deref_666_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_666_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_666_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_675_addr_0
    process(ptr_deref_675_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_675_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_675_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_675_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_675_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_675_gather_scatter
    process(ptr_deref_675_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_675_data_0;
      ov(31 downto 0) := iv;
      iNsTr_24_676 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_675_root_address_inst
    process(ptr_deref_675_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_675_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_675_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_684_addr_0
    process(ptr_deref_684_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_684_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_684_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_684_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_684_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_684_gather_scatter
    process(iNsTr_25_682) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_682;
      ov(31 downto 0) := iv;
      ptr_deref_684_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_684_root_address_inst
    process(ptr_deref_684_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_684_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_684_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_690_addr_0
    process(ptr_deref_690_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_690_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_690_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_690_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_690_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_690_gather_scatter
    process(type_cast_692_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_692_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_690_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_690_root_address_inst
    process(ptr_deref_690_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_690_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_690_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_addr_0
    process(ptr_deref_698_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_698_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_698_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_698_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_gather_scatter
    process(ptr_deref_698_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_698_data_0;
      ov(31 downto 0) := iv;
      iNsTr_28_699 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_698_root_address_inst
    process(ptr_deref_698_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_698_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_698_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_723_addr_0
    process(ptr_deref_723_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_723_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_723_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_723_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_723_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_723_gather_scatter
    process(ptr_deref_723_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_723_data_0;
      ov(31 downto 0) := iv;
      iNsTr_34_724 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_723_root_address_inst
    process(ptr_deref_723_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_723_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_723_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_737_addr_0
    process(ptr_deref_737_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_737_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_737_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_737_base_resize
    process(iNsTr_36_734) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_734;
      ov := iv(9 downto 0);
      ptr_deref_737_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_737_gather_scatter
    process(ptr_deref_737_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_737_data_0;
      ov(31 downto 0) := iv;
      iNsTr_37_738 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_737_root_address_inst
    process(ptr_deref_737_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_737_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_737_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_740_addr_0
    process(ptr_deref_740_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_740_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_740_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_740_base_resize
    process(val1_587) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val1_587;
      ov := iv(0 downto 0);
      ptr_deref_740_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_740_gather_scatter
    process(iNsTr_37_738) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_738;
      ov(31 downto 0) := iv;
      ptr_deref_740_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_740_root_address_inst
    process(ptr_deref_740_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_740_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_740_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_745_addr_0
    process(ptr_deref_745_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_745_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_745_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_745_base_resize
    process(val1_587) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val1_587;
      ov := iv(0 downto 0);
      ptr_deref_745_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_745_gather_scatter
    process(ptr_deref_745_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_745_data_0;
      ov(31 downto 0) := iv;
      iNsTr_39_746 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_745_root_address_inst
    process(ptr_deref_745_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_745_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_745_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_754_addr_0
    process(ptr_deref_754_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_754_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_754_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_754_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_754_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_754_gather_scatter
    process(ptr_deref_754_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_754_data_0;
      ov(31 downto 0) := iv;
      iNsTr_45_755 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_754_root_address_inst
    process(ptr_deref_754_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_754_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_754_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_763_addr_0
    process(ptr_deref_763_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_763_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_763_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_763_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_763_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_763_gather_scatter
    process(iNsTr_46_761) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_761;
      ov(31 downto 0) := iv;
      ptr_deref_763_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_763_root_address_inst
    process(ptr_deref_763_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_763_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_763_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_addr_0
    process(ptr_deref_769_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_769_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_769_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_769_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_gather_scatter
    process(type_cast_771_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_771_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_769_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_root_address_inst
    process(ptr_deref_769_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_769_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_769_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_777_addr_0
    process(ptr_deref_777_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_777_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_777_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_777_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_777_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_777_gather_scatter
    process(ptr_deref_777_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_777_data_0;
      ov(31 downto 0) := iv;
      iNsTr_49_778 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_777_root_address_inst
    process(ptr_deref_777_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_777_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_777_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_addr_0
    process(ptr_deref_802_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_802_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_802_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_802_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_gather_scatter
    process(ptr_deref_802_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_802_data_0;
      ov(31 downto 0) := iv;
      iNsTr_55_803 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_802_root_address_inst
    process(ptr_deref_802_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_802_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_802_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_816_addr_0
    process(ptr_deref_816_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_816_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_816_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_816_base_resize
    process(iNsTr_57_813) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_57_813;
      ov := iv(9 downto 0);
      ptr_deref_816_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_816_gather_scatter
    process(ptr_deref_816_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_816_data_0;
      ov(31 downto 0) := iv;
      iNsTr_58_817 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_816_root_address_inst
    process(ptr_deref_816_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_816_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_816_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_addr_0
    process(ptr_deref_819_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_819_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_819_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_base_resize
    process(val2_591) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val2_591;
      ov := iv(0 downto 0);
      ptr_deref_819_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_gather_scatter
    process(iNsTr_58_817) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_58_817;
      ov(31 downto 0) := iv;
      ptr_deref_819_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_root_address_inst
    process(ptr_deref_819_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_819_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_819_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_addr_0
    process(ptr_deref_824_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_824_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_824_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_base_resize
    process(val2_591) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val2_591;
      ov := iv(0 downto 0);
      ptr_deref_824_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_gather_scatter
    process(ptr_deref_824_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_824_data_0;
      ov(31 downto 0) := iv;
      iNsTr_60_825 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_824_root_address_inst
    process(ptr_deref_824_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_824_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_824_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_833_addr_0
    process(ptr_deref_833_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_833_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_833_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_833_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_833_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_833_gather_scatter
    process(ptr_deref_833_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_833_data_0;
      ov(31 downto 0) := iv;
      iNsTr_66_834 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_833_root_address_inst
    process(ptr_deref_833_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_833_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_833_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_842_addr_0
    process(ptr_deref_842_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_842_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_842_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_842_base_resize
    process(J_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_579;
      ov := iv(0 downto 0);
      ptr_deref_842_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_842_gather_scatter
    process(iNsTr_67_840) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_67_840;
      ov(31 downto 0) := iv;
      ptr_deref_842_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_842_root_address_inst
    process(ptr_deref_842_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_842_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_842_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_849_addr_0
    process(ptr_deref_849_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_849_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_849_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_849_base_resize
    process(iNsTr_0_575) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_575;
      ov := iv(0 downto 0);
      ptr_deref_849_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_849_gather_scatter
    process(ptr_deref_849_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_849_data_0;
      ov(31 downto 0) := iv;
      ret_val_x_x_buffer <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_849_root_address_inst
    process(ptr_deref_849_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_849_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_849_root_address <= ov(0 downto 0);
      --
    end process;
    if_stmt_635_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_10_634;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_635_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_635_branch_req_0,
          ack0 => if_stmt_635_branch_ack_0,
          ack1 => if_stmt_635_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_714_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_31_713;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_714_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_714_branch_req_0,
          ack0 => if_stmt_714_branch_ack_0,
          ack1 => if_stmt_714_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_793_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_52_792;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_793_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_793_branch_req_0,
          ack0 => if_stmt_793_branch_ack_0,
          ack1 => if_stmt_793_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_620_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_5_609 & iNsTr_7_616;
      iNsTr_8_621 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_620_inst_req_0;
      ADD_u32_u32_620_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_620_inst_req_1;
      ADD_u32_u32_620_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u32_u32_626_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_8_621;
      iNsTr_9_627 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_626_inst_req_0;
      ADD_u32_u32_626_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_626_inst_req_1;
      ADD_u32_u32_626_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u32_u32_681_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_24_676;
      iNsTr_25_682 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_681_inst_req_0;
      ADD_u32_u32_681_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_681_inst_req_1;
      ADD_u32_u32_681_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u32_u32_760_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_45_755;
      iNsTr_46_761 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_760_inst_req_0;
      ADD_u32_u32_760_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_760_inst_req_1;
      ADD_u32_u32_760_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ADD_u32_u32_839_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_834;
      iNsTr_67_840 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_839_inst_req_0;
      ADD_u32_u32_839_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_839_inst_req_1;
      ADD_u32_u32_839_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : SLT_i32_u1_633_inst 
    ApIntSlt_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_630_wire & type_cast_632_wire;
      iNsTr_10_634 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_633_inst_req_0;
      SLT_i32_u1_633_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_633_inst_req_1;
      SLT_i32_u1_633_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_5_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : SLT_i32_u1_712_inst 
    ApIntSlt_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_709_wire & type_cast_711_wire;
      iNsTr_31_713 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_712_inst_req_0;
      SLT_i32_u1_712_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_712_inst_req_1;
      SLT_i32_u1_712_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_6_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : SLT_i32_u1_791_inst 
    ApIntSlt_group_7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_788_wire & type_cast_790_wire;
      iNsTr_52_792 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_791_inst_req_0;
      SLT_i32_u1_791_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_791_inst_req_1;
      SLT_i32_u1_791_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_7_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : type_cast_648_inst 
    ApIntToApIntSigned_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_13_645;
      type_cast_648_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_648_inst_req_0;
      type_cast_648_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_648_inst_req_1;
      type_cast_648_inst_ack_1 <= ackR_unguarded(0);
      ApIntToApIntSigned_group_8_gI: SplitGuardInterface generic map(name => "ApIntToApIntSigned_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : type_cast_727_inst 
    ApIntToApIntSigned_group_9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_34_724;
      type_cast_727_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1 <= ackR_unguarded(0);
      ApIntToApIntSigned_group_9_gI: SplitGuardInterface generic map(name => "ApIntToApIntSigned_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : type_cast_806_inst 
    ApIntToApIntSigned_group_10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_55_803;
      type_cast_806_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_806_inst_req_0;
      type_cast_806_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_806_inst_req_1;
      type_cast_806_inst_ack_1 <= ackR_unguarded(0);
      ApIntToApIntSigned_group_10_gI: SplitGuardInterface generic map(name => "ApIntToApIntSigned_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntToApIntSigned",
          name => "ApIntToApIntSigned_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared load operator group (0) : LOAD_ncol_ind_611_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_ncol_ind_611_load_0_req_0;
      LOAD_ncol_ind_611_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ncol_ind_611_load_0_req_1;
      LOAD_ncol_ind_611_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncol_ind_611_word_address_0;
      LOAD_ncol_ind_611_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(15 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_ncols_701_load_0 LOAD_ncols_780_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= LOAD_ncols_701_load_0_req_0;
      reqL_unguarded(0) <= LOAD_ncols_780_load_0_req_0;
      LOAD_ncols_701_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_ncols_780_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_ncols_701_load_0_req_1;
      reqR_unguarded(0) <= LOAD_ncols_780_load_0_req_1;
      LOAD_ncols_701_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_ncols_780_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncols_701_word_address_0 & LOAD_ncols_780_word_address_0;
      LOAD_ncols_701_data_0 <= data_out(31 downto 16);
      LOAD_ncols_780_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_nrows_604_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_nrows_604_load_0_req_0;
      LOAD_nrows_604_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_nrows_604_load_0_req_1;
      LOAD_nrows_604_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_nrows_604_word_address_0;
      LOAD_nrows_604_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_833_load_0 ptr_deref_601_load_0 ptr_deref_644_load_0 ptr_deref_675_load_0 ptr_deref_698_load_0 ptr_deref_723_load_0 ptr_deref_754_load_0 ptr_deref_777_load_0 ptr_deref_802_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(287 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 8 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 8 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 8 downto 0);
      signal guard_vector : std_logic_vector( 8 downto 0);
      constant inBUFs : IntegerArray(8 downto 0) := (8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(8 downto 0) := (8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(8 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false);
      constant guardBuffering: IntegerArray(8 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2);
      -- 
    begin -- 
      reqL_unguarded(8) <= ptr_deref_833_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_601_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_644_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_675_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_698_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_723_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_754_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_777_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_802_load_0_req_0;
      ptr_deref_833_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_601_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_644_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_675_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_698_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_723_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_754_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_777_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_802_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(8) <= ptr_deref_833_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_601_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_644_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_675_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_698_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_723_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_754_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_777_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_802_load_0_req_1;
      ptr_deref_833_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_601_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_644_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_675_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_698_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_723_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_754_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_777_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_802_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 9, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_833_word_address_0 & ptr_deref_601_word_address_0 & ptr_deref_644_word_address_0 & ptr_deref_675_word_address_0 & ptr_deref_698_word_address_0 & ptr_deref_723_word_address_0 & ptr_deref_754_word_address_0 & ptr_deref_777_word_address_0 & ptr_deref_802_word_address_0;
      ptr_deref_833_data_0 <= data_out(287 downto 256);
      ptr_deref_601_data_0 <= data_out(255 downto 224);
      ptr_deref_644_data_0 <= data_out(223 downto 192);
      ptr_deref_675_data_0 <= data_out(191 downto 160);
      ptr_deref_698_data_0 <= data_out(159 downto 128);
      ptr_deref_723_data_0 <= data_out(127 downto 96);
      ptr_deref_754_data_0 <= data_out(95 downto 64);
      ptr_deref_777_data_0 <= data_out(63 downto 32);
      ptr_deref_802_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 9,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_19_lr_req(0),
          mack => memory_space_19_lr_ack(0),
          maddr => memory_space_19_lr_addr(0 downto 0),
          mtag => memory_space_19_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 9,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_19_lc_req(0),
          mack => memory_space_19_lc_ack(0),
          mdata => memory_space_19_lc_data(31 downto 0),
          mtag => memory_space_19_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_658_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_658_load_0_req_0;
      ptr_deref_658_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_658_load_0_req_1;
      ptr_deref_658_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_658_word_address_0;
      ptr_deref_658_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 10,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(9 downto 0),
          mtag => memory_space_4_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(15 downto 0),
          mtag => memory_space_4_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_666_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_666_load_0_req_0;
      ptr_deref_666_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_666_load_0_req_1;
      ptr_deref_666_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_666_word_address_0;
      ptr_deref_666_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_20_lr_req(0),
          mack => memory_space_20_lr_ack(0),
          maddr => memory_space_20_lr_addr(0 downto 0),
          mtag => memory_space_20_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_20_lc_req(0),
          mack => memory_space_20_lc_ack(0),
          mdata => memory_space_20_lc_data(15 downto 0),
          mtag => memory_space_20_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_737_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_737_load_0_req_0;
      ptr_deref_737_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_737_load_0_req_1;
      ptr_deref_737_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_737_word_address_0;
      ptr_deref_737_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 10,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(9 downto 0),
          mtag => memory_space_1_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_745_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_745_load_0_req_0;
      ptr_deref_745_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_745_load_0_req_1;
      ptr_deref_745_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup7_gI: SplitGuardInterface generic map(name => "LoadGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_745_word_address_0;
      ptr_deref_745_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup7", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_21_lr_req(0),
          mack => memory_space_21_lr_ack(0),
          maddr => memory_space_21_lr_addr(0 downto 0),
          mtag => memory_space_21_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup7 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_21_lc_req(0),
          mack => memory_space_21_lc_ack(0),
          mdata => memory_space_21_lc_data(31 downto 0),
          mtag => memory_space_21_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : ptr_deref_816_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_816_load_0_req_0;
      ptr_deref_816_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_816_load_0_req_1;
      ptr_deref_816_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup8_gI: SplitGuardInterface generic map(name => "LoadGroup8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_816_word_address_0;
      ptr_deref_816_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup8", addr_width => 10,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(9 downto 0),
          mtag => memory_space_0_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup8 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : ptr_deref_824_load_0 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_824_load_0_req_0;
      ptr_deref_824_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_824_load_0_req_1;
      ptr_deref_824_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup9_gI: SplitGuardInterface generic map(name => "LoadGroup9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_824_word_address_0;
      ptr_deref_824_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup9", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_22_lr_req(0),
          mack => memory_space_22_lr_ack(0),
          maddr => memory_space_22_lr_addr(0 downto 0),
          mtag => memory_space_22_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup9 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_22_lc_req(0),
          mack => memory_space_22_lc_ack(0),
          mdata => memory_space_22_lc_data(31 downto 0),
          mtag => memory_space_22_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared load operator group (10) : ptr_deref_849_load_0 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_849_load_0_req_0;
      ptr_deref_849_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_849_load_0_req_1;
      ptr_deref_849_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup10_gI: SplitGuardInterface generic map(name => "LoadGroup10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_849_word_address_0;
      ptr_deref_849_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup10", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_18_lr_req(0),
          mack => memory_space_18_lr_ack(0),
          maddr => memory_space_18_lr_addr(0 downto 0),
          mtag => memory_space_18_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup10 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_18_lc_req(0),
          mack => memory_space_18_lc_ack(0),
          mdata => memory_space_18_lc_data(31 downto 0),
          mtag => memory_space_18_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    -- shared store operator group (0) : ptr_deref_842_store_0 ptr_deref_593_store_0 ptr_deref_684_store_0 ptr_deref_690_store_0 ptr_deref_763_store_0 ptr_deref_769_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_842_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_593_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_684_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_690_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_763_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_769_store_0_req_0;
      ptr_deref_842_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_593_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_684_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_690_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_763_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_769_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_842_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_593_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_684_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_690_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_763_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_769_store_0_req_1;
      ptr_deref_842_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_593_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_684_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_690_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_763_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_769_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_842_word_address_0 & ptr_deref_593_word_address_0 & ptr_deref_684_word_address_0 & ptr_deref_690_word_address_0 & ptr_deref_763_word_address_0 & ptr_deref_769_word_address_0;
      data_in <= ptr_deref_842_data_0 & ptr_deref_593_data_0 & ptr_deref_684_data_0 & ptr_deref_690_data_0 & ptr_deref_763_data_0 & ptr_deref_769_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 6,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_19_sr_req(0),
          mack => memory_space_19_sr_ack(0),
          maddr => memory_space_19_sr_addr(0 downto 0),
          mdata => memory_space_19_sr_data(31 downto 0),
          mtag => memory_space_19_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_19_sc_req(0),
          mack => memory_space_19_sc_ack(0),
          mtag => memory_space_19_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_661_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_661_store_0_req_0;
      ptr_deref_661_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_661_store_0_req_1;
      ptr_deref_661_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_661_word_address_0;
      data_in <= ptr_deref_661_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_20_sr_req(0),
          mack => memory_space_20_sr_ack(0),
          maddr => memory_space_20_sr_addr(0 downto 0),
          mdata => memory_space_20_sr_data(15 downto 0),
          mtag => memory_space_20_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_20_sc_req(0),
          mack => memory_space_20_sc_ack(0),
          mtag => memory_space_20_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_740_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_740_store_0_req_0;
      ptr_deref_740_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_740_store_0_req_1;
      ptr_deref_740_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_740_word_address_0;
      data_in <= ptr_deref_740_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_21_sr_req(0),
          mack => memory_space_21_sr_ack(0),
          maddr => memory_space_21_sr_addr(0 downto 0),
          mdata => memory_space_21_sr_data(31 downto 0),
          mtag => memory_space_21_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_21_sc_req(0),
          mack => memory_space_21_sc_ack(0),
          mtag => memory_space_21_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_819_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_819_store_0_req_0;
      ptr_deref_819_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_819_store_0_req_1;
      ptr_deref_819_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_819_word_address_0;
      data_in <= ptr_deref_819_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_22_sr_req(0),
          mack => memory_space_22_sr_ack(0),
          maddr => memory_space_22_sr_addr(0 downto 0),
          mdata => memory_space_22_sr_data(31 downto 0),
          mtag => memory_space_22_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_22_sc_req(0),
          mack => memory_space_22_sc_ack(0),
          mtag => memory_space_22_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared outport operator group (0) : WPIPE_aPriori_out_826_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_aPriori_out_826_inst_req_0;
      WPIPE_aPriori_out_826_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_aPriori_out_826_inst_req_1;
      WPIPE_aPriori_out_826_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= iNsTr_60_825;
      aPriori_out_write_0_gI: SplitGuardInterface generic map(name => "aPriori_out_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      aPriori_out_write_0: OutputPortRevised -- 
        generic map ( name => "aPriori_out", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => aPriori_out_pipe_write_req(0),
          oack => aPriori_out_pipe_write_ack(0),
          odata => aPriori_out_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_code_block_out_747_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_code_block_out_747_inst_req_0;
      WPIPE_code_block_out_747_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_code_block_out_747_inst_req_1;
      WPIPE_code_block_out_747_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= iNsTr_39_746;
      code_block_out_write_1_gI: SplitGuardInterface generic map(name => "code_block_out_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      code_block_out_write_1: OutputPortRevised -- 
        generic map ( name => "code_block_out", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => code_block_out_pipe_write_req(0),
          oack => code_block_out_pipe_write_ack(0),
          odata => code_block_out_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_mem_out_668_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_mem_out_668_inst_req_0;
      WPIPE_mem_out_668_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_mem_out_668_inst_req_1;
      WPIPE_mem_out_668_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= iNsTr_18_667;
      mem_out_write_2_gI: SplitGuardInterface generic map(name => "mem_out_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      mem_out_write_2: OutputPortRevised -- 
        generic map ( name => "mem_out", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => mem_out_pipe_write_req(0),
          oack => mem_out_pipe_write_ack(0),
          odata => mem_out_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  dummyROM_memory_space_18: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_18",
      num_loads => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_18_lr_addr,
      lr_req_in => memory_space_18_lr_req,
      lr_ack_out => memory_space_18_lr_ack,
      lr_tag_in => memory_space_18_lr_tag,
      lc_req_in => memory_space_18_lc_req,
      lc_ack_out => memory_space_18_lc_ack,
      lc_data_out => memory_space_18_lc_data,
      lc_tag_out => memory_space_18_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_19: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_19",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_19_lr_addr,
      lr_req_in => memory_space_19_lr_req,
      lr_ack_out => memory_space_19_lr_ack,
      lr_tag_in => memory_space_19_lr_tag,
      lc_req_in => memory_space_19_lc_req,
      lc_ack_out => memory_space_19_lc_ack,
      lc_data_out => memory_space_19_lc_data,
      lc_tag_out => memory_space_19_lc_tag,
      sr_addr_in => memory_space_19_sr_addr,
      sr_data_in => memory_space_19_sr_data,
      sr_req_in => memory_space_19_sr_req,
      sr_ack_out => memory_space_19_sr_ack,
      sr_tag_in => memory_space_19_sr_tag,
      sc_req_in=> memory_space_19_sc_req,
      sc_ack_out => memory_space_19_sc_ack,
      sc_tag_out => memory_space_19_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_20: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_20",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_20_lr_addr,
      lr_req_in => memory_space_20_lr_req,
      lr_ack_out => memory_space_20_lr_ack,
      lr_tag_in => memory_space_20_lr_tag,
      lc_req_in => memory_space_20_lc_req,
      lc_ack_out => memory_space_20_lc_ack,
      lc_data_out => memory_space_20_lc_data,
      lc_tag_out => memory_space_20_lc_tag,
      sr_addr_in => memory_space_20_sr_addr,
      sr_data_in => memory_space_20_sr_data,
      sr_req_in => memory_space_20_sr_req,
      sr_ack_out => memory_space_20_sr_ack,
      sr_tag_in => memory_space_20_sr_tag,
      sc_req_in=> memory_space_20_sc_req,
      sc_ack_out => memory_space_20_sc_ack,
      sc_tag_out => memory_space_20_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_21: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_21",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_21_lr_addr,
      lr_req_in => memory_space_21_lr_req,
      lr_ack_out => memory_space_21_lr_ack,
      lr_tag_in => memory_space_21_lr_tag,
      lc_req_in => memory_space_21_lc_req,
      lc_ack_out => memory_space_21_lc_ack,
      lc_data_out => memory_space_21_lc_data,
      lc_tag_out => memory_space_21_lc_tag,
      sr_addr_in => memory_space_21_sr_addr,
      sr_data_in => memory_space_21_sr_data,
      sr_req_in => memory_space_21_sr_req,
      sr_ack_out => memory_space_21_sr_ack,
      sr_tag_in => memory_space_21_sr_tag,
      sc_req_in=> memory_space_21_sc_req,
      sc_ack_out => memory_space_21_sc_ack,
      sc_tag_out => memory_space_21_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_22: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_22",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_22_lr_addr,
      lr_req_in => memory_space_22_lr_req,
      lr_ack_out => memory_space_22_lr_ack,
      lr_tag_in => memory_space_22_lr_tag,
      lc_req_in => memory_space_22_lc_req,
      lc_ack_out => memory_space_22_lc_ack,
      lc_data_out => memory_space_22_lc_data,
      lc_tag_out => memory_space_22_lc_tag,
      sr_addr_in => memory_space_22_sr_addr,
      sr_data_in => memory_space_22_sr_data,
      sr_req_in => memory_space_22_sr_req,
      sr_ack_out => memory_space_22_sr_ack,
      sr_tag_in => memory_space_22_sr_tag,
      sc_req_in=> memory_space_22_sc_req,
      sc_ack_out => memory_space_22_sc_ack,
      sc_tag_out => memory_space_22_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end send_output_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity top_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    initInputs_call_reqs : out  std_logic_vector(0 downto 0);
    initInputs_call_acks : in   std_logic_vector(0 downto 0);
    initInputs_call_tag  :  out  std_logic_vector(0 downto 0);
    initInputs_return_reqs : out  std_logic_vector(0 downto 0);
    initInputs_return_acks : in   std_logic_vector(0 downto 0);
    initInputs_return_tag :  in   std_logic_vector(0 downto 0);
    initialize_aPriori_call_reqs : out  std_logic_vector(0 downto 0);
    initialize_aPriori_call_acks : in   std_logic_vector(0 downto 0);
    initialize_aPriori_call_tag  :  out  std_logic_vector(0 downto 0);
    initialize_aPriori_return_reqs : out  std_logic_vector(0 downto 0);
    initialize_aPriori_return_acks : in   std_logic_vector(0 downto 0);
    initialize_aPriori_return_tag :  in   std_logic_vector(0 downto 0);
    readCodeBlock_call_reqs : out  std_logic_vector(0 downto 0);
    readCodeBlock_call_acks : in   std_logic_vector(0 downto 0);
    readCodeBlock_call_tag  :  out  std_logic_vector(0 downto 0);
    readCodeBlock_return_reqs : out  std_logic_vector(0 downto 0);
    readCodeBlock_return_acks : in   std_logic_vector(0 downto 0);
    readCodeBlock_return_tag :  in   std_logic_vector(0 downto 0);
    send_output_call_reqs : out  std_logic_vector(0 downto 0);
    send_output_call_acks : in   std_logic_vector(0 downto 0);
    send_output_call_tag  :  out  std_logic_vector(0 downto 0);
    send_output_return_reqs : out  std_logic_vector(0 downto 0);
    send_output_return_acks : in   std_logic_vector(0 downto 0);
    send_output_return_data : in   std_logic_vector(31 downto 0);
    send_output_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity top_daemon;
architecture top_daemon_arch of top_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal top_daemon_CP_5761_start: Boolean;
  signal top_daemon_CP_5761_symbol: Boolean;
  -- volatile/operator module components. 
  component initInputs is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      matrix_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      matrix_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      matrix_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component initialize_aPriori is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component readCodeBlock is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      code_block_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      code_block_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      code_block_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component send_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      code_block_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      code_block_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      code_block_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      mem_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      mem_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mem_out_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_865_call_ack_1 : boolean;
  signal call_stmt_871_call_req_1 : boolean;
  signal call_stmt_871_call_ack_1 : boolean;
  signal call_stmt_871_call_req_0 : boolean;
  signal call_stmt_873_call_req_0 : boolean;
  signal call_stmt_871_call_ack_0 : boolean;
  signal ptr_deref_867_store_0_req_1 : boolean;
  signal ptr_deref_867_store_0_ack_1 : boolean;
  signal call_stmt_873_call_ack_0 : boolean;
  signal call_stmt_865_call_req_0 : boolean;
  signal call_stmt_865_call_ack_0 : boolean;
  signal call_stmt_873_call_req_1 : boolean;
  signal call_stmt_873_call_ack_1 : boolean;
  signal ptr_deref_867_store_0_req_0 : boolean;
  signal call_stmt_865_call_req_1 : boolean;
  signal ptr_deref_867_store_0_ack_0 : boolean;
  signal call_stmt_864_call_req_0 : boolean;
  signal call_stmt_864_call_ack_0 : boolean;
  signal call_stmt_864_call_req_1 : boolean;
  signal call_stmt_864_call_ack_1 : boolean;
  signal memory_space_23_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_23_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_23_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_23_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_23_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_23_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_23_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_23_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "top_daemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  top_daemon_CP_5761_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "top_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= top_daemon_CP_5761_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= top_daemon_CP_5761_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= top_daemon_CP_5761_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  top_daemon_CP_5761: Block -- control-path 
    signal top_daemon_CP_5761_elements: BooleanArray(34 downto 0);
    -- 
  begin -- 
    top_daemon_CP_5761_elements(0) <= top_daemon_CP_5761_start;
    top_daemon_CP_5761_symbol <= top_daemon_CP_5761_elements(34);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_856/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_856/branch_block_stmt_856__entry__
      -- CP-element group 1: 	 branch_block_stmt_856/assign_stmt_861__entry__
      -- 
    top_daemon_CP_5761_elements(1) <= top_daemon_CP_5761_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	27 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_856/assign_stmt_861__exit__
      -- CP-element group 2: 	 branch_block_stmt_856/bb_0_bb_1
      -- 
    top_daemon_CP_5761_elements(2) <= top_daemon_CP_5761_elements(11);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	30 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	12 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_856/merge_stmt_863__exit__
      -- CP-element group 3: 	 branch_block_stmt_856/call_stmt_864__entry__
      -- 
    top_daemon_CP_5761_elements(3) <= top_daemon_CP_5761_elements(30);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	14 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	15 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_856/call_stmt_864__exit__
      -- CP-element group 4: 	 branch_block_stmt_856/call_stmt_865__entry__
      -- 
    top_daemon_CP_5761_elements(4) <= top_daemon_CP_5761_elements(14);
    -- CP-element group 5:  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	17 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	18 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_856/call_stmt_865__exit__
      -- CP-element group 5: 	 branch_block_stmt_856/assign_stmt_870__entry__
      -- 
    top_daemon_CP_5761_elements(5) <= top_daemon_CP_5761_elements(17);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	20 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_856/assign_stmt_870__exit__
      -- CP-element group 6: 	 branch_block_stmt_856/call_stmt_871__entry__
      -- 
    top_daemon_CP_5761_elements(6) <= top_daemon_CP_5761_elements(20);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	23 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	24 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_856/call_stmt_871__exit__
      -- CP-element group 7: 	 branch_block_stmt_856/call_stmt_873__entry__
      -- 
    top_daemon_CP_5761_elements(7) <= top_daemon_CP_5761_elements(23);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	26 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	28 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_856/call_stmt_873__exit__
      -- CP-element group 8: 	 branch_block_stmt_856/bb_1_bb_1
      -- 
    top_daemon_CP_5761_elements(8) <= top_daemon_CP_5761_elements(26);
    -- CP-element group 9:  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_856/return__
      -- 
    top_daemon_CP_5761_elements(9) <= false; 
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	33 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	34 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_856/branch_block_stmt_856__exit__
      -- CP-element group 10: 	 branch_block_stmt_856/merge_stmt_876__exit__
      -- 
    top_daemon_CP_5761_elements(10) <= top_daemon_CP_5761_elements(33);
    -- CP-element group 11:  transition  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	2 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_856/assign_stmt_861/$entry
      -- CP-element group 11: 	 branch_block_stmt_856/assign_stmt_861/$exit
      -- 
    top_daemon_CP_5761_elements(11) <= top_daemon_CP_5761_elements(1);
    -- CP-element group 12:  fork  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (7) 
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/$entry
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_update_start_
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Sample/crr
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Update/ccr
      -- 
    crr_5799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(12), ack => call_stmt_864_call_req_0); -- 
    ccr_5804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(12), ack => call_stmt_864_call_req_1); -- 
    top_daemon_CP_5761_elements(12) <= top_daemon_CP_5761_elements(3);
    -- CP-element group 13:  transition  input  no-bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Sample/cra
      -- 
    cra_5800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_864_call_ack_0, ack => top_daemon_CP_5761_elements(13)); -- 
    -- CP-element group 14:  transition  input  no-bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	4 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_856/call_stmt_864/$exit
      -- CP-element group 14: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_856/call_stmt_864/call_stmt_864_Update/cca
      -- 
    cca_5805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_864_call_ack_1, ack => top_daemon_CP_5761_elements(14)); -- 
    -- CP-element group 15:  fork  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	4 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (7) 
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/$entry
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_update_start_
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Sample/crr
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Update/ccr
      -- 
    crr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(15), ack => call_stmt_865_call_req_0); -- 
    ccr_5821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(15), ack => call_stmt_865_call_req_1); -- 
    top_daemon_CP_5761_elements(15) <= top_daemon_CP_5761_elements(4);
    -- CP-element group 16:  transition  input  no-bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Sample/cra
      -- 
    cra_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_865_call_ack_0, ack => top_daemon_CP_5761_elements(16)); -- 
    -- CP-element group 17:  transition  input  no-bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	5 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Update/cca
      -- CP-element group 17: 	 branch_block_stmt_856/call_stmt_865/$exit
      -- CP-element group 17: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_856/call_stmt_865/call_stmt_865_Update/$exit
      -- 
    cca_5822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_865_call_ack_1, ack => top_daemon_CP_5761_elements(17)); -- 
    -- CP-element group 18:  join  fork  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	5 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (31) 
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_update_start_
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/word_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/ptr_deref_867_Split/split_ack
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_address_resized
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/ptr_deref_867_Split/split_req
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_addr_resize/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/word_0/cr
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_addr_resize/$exit
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_addr_resize/base_resize_req
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_addr_resize/base_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/ptr_deref_867_Split/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/word_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/ptr_deref_867_Split/$exit
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/word_0/rr
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_word_addrgen/$entry
      -- 
    cr_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(18), ack => ptr_deref_867_store_0_req_1); -- 
    rr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(18), ack => ptr_deref_867_store_0_req_0); -- 
    top_daemon_CP_5761_elements(18) <= top_daemon_CP_5761_elements(5);
    -- CP-element group 19:  transition  input  no-bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Sample/word_access_start/word_0/ra
      -- 
    ra_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_867_store_0_ack_0, ack => top_daemon_CP_5761_elements(19)); -- 
    -- CP-element group 20:  transition  input  no-bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	6 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/$exit
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_856/assign_stmt_870/ptr_deref_867_Update/word_access_complete/word_0/ca
      -- 
    ca_5875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_867_store_0_ack_1, ack => top_daemon_CP_5761_elements(20)); -- 
    -- CP-element group 21:  fork  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (7) 
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Update/ccr
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Sample/crr
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/$entry
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_update_start_
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_sample_start_
      -- 
    crr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(21), ack => call_stmt_871_call_req_0); -- 
    ccr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(21), ack => call_stmt_871_call_req_1); -- 
    top_daemon_CP_5761_elements(21) <= top_daemon_CP_5761_elements(6);
    -- CP-element group 22:  transition  input  no-bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Sample/cra
      -- 
    cra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_871_call_ack_0, ack => top_daemon_CP_5761_elements(22)); -- 
    -- CP-element group 23:  transition  input  no-bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	7 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_Update/cca
      -- CP-element group 23: 	 branch_block_stmt_856/call_stmt_871/$exit
      -- CP-element group 23: 	 branch_block_stmt_856/call_stmt_871/call_stmt_871_update_completed_
      -- 
    cca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_871_call_ack_1, ack => top_daemon_CP_5761_elements(23)); -- 
    -- CP-element group 24:  fork  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	7 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (7) 
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Sample/crr
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/$entry
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Update/ccr
      -- CP-element group 24: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_update_start_
      -- 
    crr_5903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(24), ack => call_stmt_873_call_req_0); -- 
    ccr_5908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => top_daemon_CP_5761_elements(24), ack => call_stmt_873_call_req_1); -- 
    top_daemon_CP_5761_elements(24) <= top_daemon_CP_5761_elements(7);
    -- CP-element group 25:  transition  input  no-bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Sample/cra
      -- 
    cra_5904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_873_call_ack_0, ack => top_daemon_CP_5761_elements(25)); -- 
    -- CP-element group 26:  transition  input  no-bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	8 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_856/call_stmt_873/$exit
      -- CP-element group 26: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_856/call_stmt_873/call_stmt_873_Update/cca
      -- 
    cca_5909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_873_call_ack_1, ack => top_daemon_CP_5761_elements(26)); -- 
    -- CP-element group 27:  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_856/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_856/bb_0_bb_1_PhiReq/$exit
      -- 
    top_daemon_CP_5761_elements(27) <= top_daemon_CP_5761_elements(2);
    -- CP-element group 28:  transition  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	8 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_856/bb_1_bb_1_PhiReq/$entry
      -- CP-element group 28: 	 branch_block_stmt_856/bb_1_bb_1_PhiReq/$exit
      -- 
    top_daemon_CP_5761_elements(28) <= top_daemon_CP_5761_elements(8);
    -- CP-element group 29:  merge  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_856/merge_stmt_863_PhiReqMerge
      -- 
    top_daemon_CP_5761_elements(29) <= OrReduce(top_daemon_CP_5761_elements(27) & top_daemon_CP_5761_elements(28));
    -- CP-element group 30:  transition  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	3 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_856/merge_stmt_863_PhiAck/$entry
      -- CP-element group 30: 	 branch_block_stmt_856/merge_stmt_863_PhiAck/$exit
      -- CP-element group 30: 	 branch_block_stmt_856/merge_stmt_863_PhiAck/dummy
      -- 
    top_daemon_CP_5761_elements(30) <= top_daemon_CP_5761_elements(29);
    -- CP-element group 31:  transition  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_856/return___PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_856/return___PhiReq/$exit
      -- 
    top_daemon_CP_5761_elements(31) <= top_daemon_CP_5761_elements(9);
    -- CP-element group 32:  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_856/merge_stmt_876_PhiReqMerge
      -- 
    top_daemon_CP_5761_elements(32) <= top_daemon_CP_5761_elements(31);
    -- CP-element group 33:  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	10 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_856/merge_stmt_876_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_856/merge_stmt_876_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_856/merge_stmt_876_PhiAck/dummy
      -- 
    top_daemon_CP_5761_elements(33) <= top_daemon_CP_5761_elements(32);
    -- CP-element group 34:  transition  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	10 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 $exit
      -- CP-element group 34: 	 branch_block_stmt_856/$exit
      -- 
    top_daemon_CP_5761_elements(34) <= top_daemon_CP_5761_elements(10);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal iNsTr_5_873 : std_logic_vector(31 downto 0);
    signal nitr_861 : std_logic_vector(31 downto 0);
    signal ptr_deref_867_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_867_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_867_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_867_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_867_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_867_word_offset_0 : std_logic_vector(0 downto 0);
    signal type_cast_869_wire_constant : std_logic_vector(7 downto 0);
    signal xxtop_daemonxxbodyxxnitr_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    nitr_861 <= "00000000000000000000000000000000";
    ptr_deref_867_word_offset_0 <= "0";
    type_cast_869_wire_constant <= "00000001";
    xxtop_daemonxxbodyxxnitr_alloc_base_address <= "0";
    -- equivalence ptr_deref_867_addr_0
    process(ptr_deref_867_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_867_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_867_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_867_base_resize
    process(nitr_861) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := nitr_861;
      ov := iv(0 downto 0);
      ptr_deref_867_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_867_gather_scatter
    process(type_cast_869_wire_constant) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_869_wire_constant;
      ov(7 downto 0) := iv;
      ptr_deref_867_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_867_root_address_inst
    process(ptr_deref_867_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_867_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_867_root_address <= ov(0 downto 0);
      --
    end process;
    -- shared store operator group (0) : ptr_deref_867_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_867_store_0_req_0;
      ptr_deref_867_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_867_store_0_req_1;
      ptr_deref_867_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_867_word_address_0;
      data_in <= ptr_deref_867_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_23_sr_req(0),
          mack => memory_space_23_sr_ack(0),
          maddr => memory_space_23_sr_addr(0 downto 0),
          mdata => memory_space_23_sr_data(7 downto 0),
          mtag => memory_space_23_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_23_sc_req(0),
          mack => memory_space_23_sc_ack(0),
          mtag => memory_space_23_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared call operator group (0) : call_stmt_864_call 
    initInputs_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_864_call_req_0;
      call_stmt_864_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_864_call_req_1;
      call_stmt_864_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initInputs_call_group_0_gI: SplitGuardInterface generic map(name => "initInputs_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => initInputs_call_reqs(0),
          ackR => initInputs_call_acks(0),
          tagR => initInputs_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => initInputs_return_acks(0), -- cross-over
          ackL => initInputs_return_reqs(0), -- cross-over
          tagL => initInputs_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_865_call 
    readCodeBlock_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_865_call_req_0;
      call_stmt_865_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_865_call_req_1;
      call_stmt_865_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readCodeBlock_call_group_1_gI: SplitGuardInterface generic map(name => "readCodeBlock_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => readCodeBlock_call_reqs(0),
          ackR => readCodeBlock_call_acks(0),
          tagR => readCodeBlock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => readCodeBlock_return_acks(0), -- cross-over
          ackL => readCodeBlock_return_reqs(0), -- cross-over
          tagL => readCodeBlock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_871_call 
    initialize_aPriori_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_871_call_req_0;
      call_stmt_871_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_871_call_req_1;
      call_stmt_871_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initialize_aPriori_call_group_2_gI: SplitGuardInterface generic map(name => "initialize_aPriori_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => initialize_aPriori_call_reqs(0),
          ackR => initialize_aPriori_call_acks(0),
          tagR => initialize_aPriori_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => initialize_aPriori_return_acks(0), -- cross-over
          ackL => initialize_aPriori_return_reqs(0), -- cross-over
          tagL => initialize_aPriori_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_873_call 
    send_output_call_group_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_873_call_req_0;
      call_stmt_873_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_873_call_req_1;
      call_stmt_873_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      send_output_call_group_3_gI: SplitGuardInterface generic map(name => "send_output_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      iNsTr_5_873 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => send_output_call_reqs(0),
          ackR => send_output_call_acks(0),
          tagR => send_output_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => send_output_return_acks(0), -- cross-over
          ackL => send_output_return_reqs(0), -- cross-over
          dataL => send_output_return_data(31 downto 0),
          tagL => send_output_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  dummyWOM_memory_space_23: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_23",
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_23_sr_addr,
      sr_data_in => memory_space_23_sr_data,
      sr_req_in => memory_space_23_sr_req,
      sr_ack_out => memory_space_23_sr_ack,
      sr_tag_in => memory_space_23_sr_tag,
      sc_req_in=> memory_space_23_sc_req,
      sc_ack_out => memory_space_23_sc_ack,
      sc_tag_out => memory_space_23_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end top_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    aPriori_out_pipe_read_data: out std_logic_vector(31 downto 0);
    aPriori_out_pipe_read_req : in std_logic_vector(0 downto 0);
    aPriori_out_pipe_read_ack : out std_logic_vector(0 downto 0);
    code_block_in_pipe_write_data: in std_logic_vector(31 downto 0);
    code_block_in_pipe_write_req : in std_logic_vector(0 downto 0);
    code_block_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    code_block_out_pipe_read_data: out std_logic_vector(31 downto 0);
    code_block_out_pipe_read_req : in std_logic_vector(0 downto 0);
    code_block_out_pipe_read_ack : out std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_write_data: in std_logic_vector(31 downto 0);
    ebbyNo_in_pipe_write_req : in std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    matrix_in_pipe_write_data: in std_logic_vector(15 downto 0);
    matrix_in_pipe_write_req : in std_logic_vector(0 downto 0);
    matrix_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxNitr_in_pipe_write_data: in std_logic_vector(15 downto 0);
    maxNitr_in_pipe_write_req : in std_logic_vector(0 downto 0);
    maxNitr_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    mem_out_pipe_read_data: out std_logic_vector(15 downto 0);
    mem_out_pipe_read_req : in std_logic_vector(0 downto 0);
    mem_out_pipe_read_ack : out std_logic_vector(0 downto 0);
    rate_in_pipe_write_data: in std_logic_vector(31 downto 0);
    rate_in_pipe_write_req : in std_logic_vector(0 downto 0);
    rate_in_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(19 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(11 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(47 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module initInputs
  component initInputs is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      matrix_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      matrix_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      matrix_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initInputs
  signal initInputs_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initInputs_tag_out   : std_logic_vector(1 downto 0);
  signal initInputs_start_req : std_logic;
  signal initInputs_start_ack : std_logic;
  signal initInputs_fin_req   : std_logic;
  signal initInputs_fin_ack : std_logic;
  -- caller side aggregated signals for module initInputs
  signal initInputs_call_reqs: std_logic_vector(0 downto 0);
  signal initInputs_call_acks: std_logic_vector(0 downto 0);
  signal initInputs_return_reqs: std_logic_vector(0 downto 0);
  signal initInputs_return_acks: std_logic_vector(0 downto 0);
  signal initInputs_call_tag: std_logic_vector(0 downto 0);
  signal initInputs_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module initialize_aPriori
  component initialize_aPriori is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initialize_aPriori
  signal initialize_aPriori_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initialize_aPriori_tag_out   : std_logic_vector(1 downto 0);
  signal initialize_aPriori_start_req : std_logic;
  signal initialize_aPriori_start_ack : std_logic;
  signal initialize_aPriori_fin_req   : std_logic;
  signal initialize_aPriori_fin_ack : std_logic;
  -- caller side aggregated signals for module initialize_aPriori
  signal initialize_aPriori_call_reqs: std_logic_vector(0 downto 0);
  signal initialize_aPriori_call_acks: std_logic_vector(0 downto 0);
  signal initialize_aPriori_return_reqs: std_logic_vector(0 downto 0);
  signal initialize_aPriori_return_acks: std_logic_vector(0 downto 0);
  signal initialize_aPriori_call_tag: std_logic_vector(0 downto 0);
  signal initialize_aPriori_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module readCodeBlock
  component readCodeBlock is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      code_block_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      code_block_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      code_block_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readCodeBlock
  signal readCodeBlock_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readCodeBlock_tag_out   : std_logic_vector(1 downto 0);
  signal readCodeBlock_start_req : std_logic;
  signal readCodeBlock_start_ack : std_logic;
  signal readCodeBlock_fin_req   : std_logic;
  signal readCodeBlock_fin_ack : std_logic;
  -- caller side aggregated signals for module readCodeBlock
  signal readCodeBlock_call_reqs: std_logic_vector(0 downto 0);
  signal readCodeBlock_call_acks: std_logic_vector(0 downto 0);
  signal readCodeBlock_return_reqs: std_logic_vector(0 downto 0);
  signal readCodeBlock_return_acks: std_logic_vector(0 downto 0);
  signal readCodeBlock_call_tag: std_logic_vector(0 downto 0);
  signal readCodeBlock_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module send_output
  component send_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(31 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      aPriori_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      code_block_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      code_block_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      code_block_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      mem_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      mem_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mem_out_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module send_output
  signal send_output_ret_val_x_x :  std_logic_vector(31 downto 0);
  signal send_output_out_args   : std_logic_vector(31 downto 0);
  signal send_output_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal send_output_tag_out   : std_logic_vector(1 downto 0);
  signal send_output_start_req : std_logic;
  signal send_output_start_ack : std_logic;
  signal send_output_fin_req   : std_logic;
  signal send_output_fin_ack : std_logic;
  -- caller side aggregated signals for module send_output
  signal send_output_call_reqs: std_logic_vector(0 downto 0);
  signal send_output_call_acks: std_logic_vector(0 downto 0);
  signal send_output_return_reqs: std_logic_vector(0 downto 0);
  signal send_output_return_acks: std_logic_vector(0 downto 0);
  signal send_output_call_tag: std_logic_vector(0 downto 0);
  signal send_output_return_data: std_logic_vector(31 downto 0);
  signal send_output_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module top_daemon
  component top_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      initInputs_call_reqs : out  std_logic_vector(0 downto 0);
      initInputs_call_acks : in   std_logic_vector(0 downto 0);
      initInputs_call_tag  :  out  std_logic_vector(0 downto 0);
      initInputs_return_reqs : out  std_logic_vector(0 downto 0);
      initInputs_return_acks : in   std_logic_vector(0 downto 0);
      initInputs_return_tag :  in   std_logic_vector(0 downto 0);
      initialize_aPriori_call_reqs : out  std_logic_vector(0 downto 0);
      initialize_aPriori_call_acks : in   std_logic_vector(0 downto 0);
      initialize_aPriori_call_tag  :  out  std_logic_vector(0 downto 0);
      initialize_aPriori_return_reqs : out  std_logic_vector(0 downto 0);
      initialize_aPriori_return_acks : in   std_logic_vector(0 downto 0);
      initialize_aPriori_return_tag :  in   std_logic_vector(0 downto 0);
      readCodeBlock_call_reqs : out  std_logic_vector(0 downto 0);
      readCodeBlock_call_acks : in   std_logic_vector(0 downto 0);
      readCodeBlock_call_tag  :  out  std_logic_vector(0 downto 0);
      readCodeBlock_return_reqs : out  std_logic_vector(0 downto 0);
      readCodeBlock_return_acks : in   std_logic_vector(0 downto 0);
      readCodeBlock_return_tag :  in   std_logic_vector(0 downto 0);
      send_output_call_reqs : out  std_logic_vector(0 downto 0);
      send_output_call_acks : in   std_logic_vector(0 downto 0);
      send_output_call_tag  :  out  std_logic_vector(0 downto 0);
      send_output_return_reqs : out  std_logic_vector(0 downto 0);
      send_output_return_acks : in   std_logic_vector(0 downto 0);
      send_output_return_data : in   std_logic_vector(31 downto 0);
      send_output_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module top_daemon
  signal top_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal top_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal top_daemon_start_req : std_logic;
  signal top_daemon_start_ack : std_logic;
  signal top_daemon_fin_req   : std_logic;
  signal top_daemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe aPriori_out
  signal aPriori_out_pipe_write_data: std_logic_vector(31 downto 0);
  signal aPriori_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal aPriori_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe code_block_in
  signal code_block_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal code_block_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal code_block_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe code_block_out
  signal code_block_out_pipe_write_data: std_logic_vector(31 downto 0);
  signal code_block_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal code_block_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ebbyNo_in
  signal ebbyNo_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal ebbyNo_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal ebbyNo_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe matrix_in
  signal matrix_in_pipe_read_data: std_logic_vector(15 downto 0);
  signal matrix_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal matrix_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxNitr_in
  signal maxNitr_in_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxNitr_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxNitr_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe mem_out
  signal mem_out_pipe_write_data: std_logic_vector(15 downto 0);
  signal mem_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal mem_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe rate_in
  signal rate_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal rate_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal rate_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module initInputs
  -- call arbiter for module initInputs
  initInputs_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initInputs_call_reqs,
      call_acks => initInputs_call_acks,
      return_reqs => initInputs_return_reqs,
      return_acks => initInputs_return_acks,
      call_tag  => initInputs_call_tag,
      return_tag  => initInputs_return_tag,
      call_mtag => initInputs_tag_in,
      return_mtag => initInputs_tag_out,
      call_mreq => initInputs_start_req,
      call_mack => initInputs_start_ack,
      return_mreq => initInputs_fin_req,
      return_mack => initInputs_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  initInputs_instance:initInputs-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => initInputs_start_req,
      start_ack => initInputs_start_ack,
      fin_req => initInputs_fin_req,
      fin_ack => initInputs_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(19 downto 10),
      memory_space_4_lr_tag => memory_space_4_lr_tag(11 downto 6),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 16),
      memory_space_4_lc_tag => memory_space_4_lc_tag(5 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(0 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(15 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(0 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(9 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(15 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(5 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(2 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(0 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(15 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(3 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(5 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(3 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(31 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(0 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(0 downto 0),
      ebbyNo_in_pipe_read_req => ebbyNo_in_pipe_read_req(0 downto 0),
      ebbyNo_in_pipe_read_ack => ebbyNo_in_pipe_read_ack(0 downto 0),
      ebbyNo_in_pipe_read_data => ebbyNo_in_pipe_read_data(31 downto 0),
      rate_in_pipe_read_req => rate_in_pipe_read_req(0 downto 0),
      rate_in_pipe_read_ack => rate_in_pipe_read_ack(0 downto 0),
      rate_in_pipe_read_data => rate_in_pipe_read_data(31 downto 0),
      matrix_in_pipe_read_req => matrix_in_pipe_read_req(0 downto 0),
      matrix_in_pipe_read_ack => matrix_in_pipe_read_ack(0 downto 0),
      matrix_in_pipe_read_data => matrix_in_pipe_read_data(15 downto 0),
      maxNitr_in_pipe_read_req => maxNitr_in_pipe_read_req(0 downto 0),
      maxNitr_in_pipe_read_ack => maxNitr_in_pipe_read_ack(0 downto 0),
      maxNitr_in_pipe_read_data => maxNitr_in_pipe_read_data(15 downto 0),
      tag_in => initInputs_tag_in,
      tag_out => initInputs_tag_out-- 
    ); -- 
  -- module initialize_aPriori
  -- call arbiter for module initialize_aPriori
  initialize_aPriori_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initialize_aPriori_call_reqs,
      call_acks => initialize_aPriori_call_acks,
      return_reqs => initialize_aPriori_return_reqs,
      return_acks => initialize_aPriori_return_acks,
      call_tag  => initialize_aPriori_call_tag,
      return_tag  => initialize_aPriori_return_tag,
      call_mtag => initialize_aPriori_tag_in,
      return_mtag => initialize_aPriori_tag_out,
      call_mreq => initialize_aPriori_start_req,
      call_mack => initialize_aPriori_start_ack,
      return_mreq => initialize_aPriori_fin_req,
      return_mack => initialize_aPriori_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  initialize_aPriori_instance:initialize_aPriori-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => initialize_aPriori_start_req,
      start_ack => initialize_aPriori_start_ack,
      fin_req => initialize_aPriori_fin_req,
      fin_ack => initialize_aPriori_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_6_lr_req => memory_space_6_lr_req(2 downto 2),
      memory_space_6_lr_ack => memory_space_6_lr_ack(2 downto 2),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 2),
      memory_space_6_lr_tag => memory_space_6_lr_tag(17 downto 12),
      memory_space_6_lc_req => memory_space_6_lc_req(2 downto 2),
      memory_space_6_lc_ack => memory_space_6_lc_ack(2 downto 2),
      memory_space_6_lc_data => memory_space_6_lc_data(47 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(5 downto 4),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(9 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(3 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => initialize_aPriori_tag_in,
      tag_out => initialize_aPriori_tag_out-- 
    ); -- 
  -- module readCodeBlock
  -- call arbiter for module readCodeBlock
  readCodeBlock_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readCodeBlock_call_reqs,
      call_acks => readCodeBlock_call_acks,
      return_reqs => readCodeBlock_return_reqs,
      return_acks => readCodeBlock_return_acks,
      call_tag  => readCodeBlock_call_tag,
      return_tag  => readCodeBlock_return_tag,
      call_mtag => readCodeBlock_tag_in,
      return_mtag => readCodeBlock_tag_out,
      call_mreq => readCodeBlock_start_req,
      call_mack => readCodeBlock_start_ack,
      return_mreq => readCodeBlock_fin_req,
      return_mack => readCodeBlock_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  readCodeBlock_instance:readCodeBlock-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => readCodeBlock_start_req,
      start_ack => readCodeBlock_start_ack,
      fin_req => readCodeBlock_fin_req,
      fin_ack => readCodeBlock_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(11 downto 6),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 16),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(9 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(3 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      code_block_in_pipe_read_req => code_block_in_pipe_read_req(0 downto 0),
      code_block_in_pipe_read_ack => code_block_in_pipe_read_ack(0 downto 0),
      code_block_in_pipe_read_data => code_block_in_pipe_read_data(31 downto 0),
      tag_in => readCodeBlock_tag_in,
      tag_out => readCodeBlock_tag_out-- 
    ); -- 
  -- module send_output
  send_output_out_args <= send_output_ret_val_x_x ;
  -- call arbiter for module send_output
  send_output_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => send_output_call_reqs,
      call_acks => send_output_call_acks,
      return_reqs => send_output_return_reqs,
      return_acks => send_output_return_acks,
      call_tag  => send_output_call_tag,
      return_tag  => send_output_return_tag,
      call_mtag => send_output_tag_in,
      return_mtag => send_output_tag_out,
      return_data =>send_output_return_data,
      call_mreq => send_output_start_req,
      call_mack => send_output_start_ack,
      return_mreq => send_output_fin_req,
      return_mack => send_output_fin_ack,
      return_mdata => send_output_out_args,
      clk => clk, 
      reset => reset --
    ); --
  send_output_instance:send_output-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => send_output_ret_val_x_x,
      start_req => send_output_start_req,
      start_ack => send_output_start_ack,
      fin_req => send_output_fin_req,
      fin_ack => send_output_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(9 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(3 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(9 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(3 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(9 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(5 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(15 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(0 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(3 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(15 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(5 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(3 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      aPriori_out_pipe_write_req => aPriori_out_pipe_write_req(0 downto 0),
      aPriori_out_pipe_write_ack => aPriori_out_pipe_write_ack(0 downto 0),
      aPriori_out_pipe_write_data => aPriori_out_pipe_write_data(31 downto 0),
      code_block_out_pipe_write_req => code_block_out_pipe_write_req(0 downto 0),
      code_block_out_pipe_write_ack => code_block_out_pipe_write_ack(0 downto 0),
      code_block_out_pipe_write_data => code_block_out_pipe_write_data(31 downto 0),
      mem_out_pipe_write_req => mem_out_pipe_write_req(0 downto 0),
      mem_out_pipe_write_ack => mem_out_pipe_write_ack(0 downto 0),
      mem_out_pipe_write_data => mem_out_pipe_write_data(15 downto 0),
      tag_in => send_output_tag_in,
      tag_out => send_output_tag_out-- 
    ); -- 
  -- module top_daemon
  top_daemon_instance:top_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => top_daemon_start_req,
      start_ack => top_daemon_start_ack,
      fin_req => top_daemon_fin_req,
      fin_ack => top_daemon_fin_ack,
      clk => clk,
      reset => reset,
      initInputs_call_reqs => initInputs_call_reqs(0 downto 0),
      initInputs_call_acks => initInputs_call_acks(0 downto 0),
      initInputs_call_tag => initInputs_call_tag(0 downto 0),
      initInputs_return_reqs => initInputs_return_reqs(0 downto 0),
      initInputs_return_acks => initInputs_return_acks(0 downto 0),
      initInputs_return_tag => initInputs_return_tag(0 downto 0),
      initialize_aPriori_call_reqs => initialize_aPriori_call_reqs(0 downto 0),
      initialize_aPriori_call_acks => initialize_aPriori_call_acks(0 downto 0),
      initialize_aPriori_call_tag => initialize_aPriori_call_tag(0 downto 0),
      initialize_aPriori_return_reqs => initialize_aPriori_return_reqs(0 downto 0),
      initialize_aPriori_return_acks => initialize_aPriori_return_acks(0 downto 0),
      initialize_aPriori_return_tag => initialize_aPriori_return_tag(0 downto 0),
      readCodeBlock_call_reqs => readCodeBlock_call_reqs(0 downto 0),
      readCodeBlock_call_acks => readCodeBlock_call_acks(0 downto 0),
      readCodeBlock_call_tag => readCodeBlock_call_tag(0 downto 0),
      readCodeBlock_return_reqs => readCodeBlock_return_reqs(0 downto 0),
      readCodeBlock_return_acks => readCodeBlock_return_acks(0 downto 0),
      readCodeBlock_return_tag => readCodeBlock_return_tag(0 downto 0),
      send_output_call_reqs => send_output_call_reqs(0 downto 0),
      send_output_call_acks => send_output_call_acks(0 downto 0),
      send_output_call_tag => send_output_call_tag(0 downto 0),
      send_output_return_reqs => send_output_return_reqs(0 downto 0),
      send_output_return_acks => send_output_return_acks(0 downto 0),
      send_output_return_data => send_output_return_data(31 downto 0),
      send_output_return_tag => send_output_return_tag(0 downto 0),
      tag_in => top_daemon_tag_in,
      tag_out => top_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  top_daemon_tag_in <= (others => '0');
  top_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => top_daemon_start_req, start_ack => top_daemon_start_ack,  fin_req => top_daemon_fin_req,  fin_ack => top_daemon_fin_ack);
  aPriori_out_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe aPriori_out",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => aPriori_out_pipe_read_req,
      read_ack => aPriori_out_pipe_read_ack,
      read_data => aPriori_out_pipe_read_data,
      write_req => aPriori_out_pipe_write_req,
      write_ack => aPriori_out_pipe_write_ack,
      write_data => aPriori_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  code_block_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe code_block_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => code_block_in_pipe_read_req,
      read_ack => code_block_in_pipe_read_ack,
      read_data => code_block_in_pipe_read_data,
      write_req => code_block_in_pipe_write_req,
      write_ack => code_block_in_pipe_write_ack,
      write_data => code_block_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  code_block_out_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe code_block_out",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => code_block_out_pipe_read_req,
      read_ack => code_block_out_pipe_read_ack,
      read_data => code_block_out_pipe_read_data,
      write_req => code_block_out_pipe_write_req,
      write_ack => code_block_out_pipe_write_ack,
      write_data => code_block_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ebbyNo_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ebbyNo_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ebbyNo_in_pipe_read_req,
      read_ack => ebbyNo_in_pipe_read_ack,
      read_data => ebbyNo_in_pipe_read_data,
      write_req => ebbyNo_in_pipe_write_req,
      write_ack => ebbyNo_in_pipe_write_ack,
      write_data => ebbyNo_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  matrix_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe matrix_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => matrix_in_pipe_read_req,
      read_ack => matrix_in_pipe_read_ack,
      read_data => matrix_in_pipe_read_data,
      write_req => matrix_in_pipe_write_req,
      write_ack => matrix_in_pipe_write_ack,
      write_data => matrix_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxNitr_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxNitr_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxNitr_in_pipe_read_req,
      read_ack => maxNitr_in_pipe_read_ack,
      read_data => maxNitr_in_pipe_read_data,
      write_req => maxNitr_in_pipe_write_req,
      write_ack => maxNitr_in_pipe_write_ack,
      write_data => maxNitr_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mem_out_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mem_out",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => mem_out_pipe_read_req,
      read_ack => mem_out_pipe_read_ack,
      read_data => mem_out_pipe_read_data,
      write_req => mem_out_pipe_write_req,
      write_ack => mem_out_pipe_write_ack,
      write_data => mem_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  rate_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe rate_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => rate_in_pipe_read_req,
      read_ack => rate_in_pipe_read_ack,
      read_data => rate_in_pipe_read_data,
      write_req => rate_in_pipe_write_req,
      write_ack => rate_in_pipe_write_ack,
      write_data => rate_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_3: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 2,
      num_stores => 1,
      addr_width => 10,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 3,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 4,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_8: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
