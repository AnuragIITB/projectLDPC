-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity checkNodeComputeEngine is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_9_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_9_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_9_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_9_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_10_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_12_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_12_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_12_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_12_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_12_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_12_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity checkNodeComputeEngine;
architecture checkNodeComputeEngine_arch of checkNodeComputeEngine is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal checkNodeComputeEngine_CP_1062_start: Boolean;
  signal checkNodeComputeEngine_CP_1062_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal EQ_u16_u1_386_inst_ack_0 : boolean;
  signal ADD_u64_u64_403_inst_ack_0 : boolean;
  signal ADD_u64_u64_403_inst_req_0 : boolean;
  signal ADD_u64_u64_326_inst_req_0 : boolean;
  signal if_stmt_680_branch_ack_1 : boolean;
  signal type_cast_397_inst_ack_1 : boolean;
  signal ADD_u64_u64_321_inst_ack_0 : boolean;
  signal ADD_u64_u64_321_inst_req_0 : boolean;
  signal SUB_u16_u16_349_inst_ack_1 : boolean;
  signal EQ_u16_u1_386_inst_req_0 : boolean;
  signal ADD_u16_u16_366_inst_ack_0 : boolean;
  signal ADD_u64_u64_303_inst_ack_0 : boolean;
  signal type_cast_397_inst_ack_0 : boolean;
  signal addr_of_356_final_reg_ack_0 : boolean;
  signal ptr_deref_344_load_0_req_0 : boolean;
  signal ptr_deref_344_load_0_ack_0 : boolean;
  signal ptr_deref_360_load_0_req_1 : boolean;
  signal ADD_u64_u64_303_inst_req_0 : boolean;
  signal ptr_deref_360_load_0_ack_1 : boolean;
  signal addr_of_331_final_reg_req_0 : boolean;
  signal EQ_u16_u1_386_inst_req_1 : boolean;
  signal ptr_deref_360_load_0_req_0 : boolean;
  signal if_stmt_310_branch_ack_1 : boolean;
  signal EQ_u16_u1_386_inst_ack_1 : boolean;
  signal if_stmt_388_branch_ack_0 : boolean;
  signal ADD_u16_u16_366_inst_ack_1 : boolean;
  signal ADD_u16_u16_366_inst_req_1 : boolean;
  signal SUB_u16_u16_349_inst_ack_0 : boolean;
  signal ADD_u64_u64_326_inst_ack_0 : boolean;
  signal ptr_deref_340_load_0_req_0 : boolean;
  signal ptr_deref_344_load_0_req_1 : boolean;
  signal addr_of_356_final_reg_req_0 : boolean;
  signal ptr_deref_340_load_0_ack_0 : boolean;
  signal ADD_u64_u64_303_inst_req_1 : boolean;
  signal ptr_deref_344_load_0_ack_1 : boolean;
  signal if_stmt_310_branch_req_0 : boolean;
  signal ptr_deref_340_load_0_req_1 : boolean;
  signal ptr_deref_340_load_0_ack_1 : boolean;
  signal addr_of_331_final_reg_ack_0 : boolean;
  signal SUB_u16_u16_371_inst_req_0 : boolean;
  signal type_cast_397_inst_req_1 : boolean;
  signal SUB_u16_u16_371_inst_ack_0 : boolean;
  signal if_stmt_388_branch_req_0 : boolean;
  signal ADD_u64_u64_303_inst_ack_1 : boolean;
  signal addr_of_356_final_reg_req_1 : boolean;
  signal addr_of_356_final_reg_ack_1 : boolean;
  signal ADD_u64_u64_308_inst_req_0 : boolean;
  signal if_stmt_388_branch_ack_1 : boolean;
  signal SUB_u16_u16_371_inst_req_1 : boolean;
  signal SUB_u16_u16_371_inst_ack_1 : boolean;
  signal ADD_u16_u16_366_inst_req_0 : boolean;
  signal if_stmt_310_branch_ack_0 : boolean;
  signal SUB_u16_u16_349_inst_req_0 : boolean;
  signal SUB_u16_u16_349_inst_req_1 : boolean;
  signal ADD_u64_u64_321_inst_req_1 : boolean;
  signal addr_of_331_final_reg_req_1 : boolean;
  signal ADD_u64_u64_308_inst_ack_0 : boolean;
  signal ADD_u64_u64_321_inst_ack_1 : boolean;
  signal addr_of_336_final_reg_req_0 : boolean;
  signal addr_of_336_final_reg_ack_0 : boolean;
  signal ptr_deref_360_load_0_ack_0 : boolean;
  signal ADD_u64_u64_308_inst_req_1 : boolean;
  signal addr_of_336_final_reg_req_1 : boolean;
  signal ADD_u64_u64_326_inst_req_1 : boolean;
  signal ADD_u64_u64_308_inst_ack_1 : boolean;
  signal addr_of_336_final_reg_ack_1 : boolean;
  signal addr_of_331_final_reg_ack_1 : boolean;
  signal type_cast_397_inst_req_0 : boolean;
  signal ADD_u64_u64_326_inst_ack_1 : boolean;
  signal ULT_u16_u1_692_inst_ack_0 : boolean;
  signal if_stmt_680_branch_ack_0 : boolean;
  signal addr_of_663_final_reg_req_0 : boolean;
  signal LOAD_nrows_228_load_0_req_0 : boolean;
  signal LOAD_nrows_228_load_0_ack_0 : boolean;
  signal LOAD_nrows_228_load_0_req_1 : boolean;
  signal LOAD_nrows_228_load_0_ack_1 : boolean;
  signal ADD_u16_u16_673_inst_req_0 : boolean;
  signal ADD_u16_u16_673_inst_ack_0 : boolean;
  signal EQ_u16_u1_234_inst_req_0 : boolean;
  signal EQ_u16_u1_234_inst_ack_0 : boolean;
  signal EQ_u16_u1_234_inst_req_1 : boolean;
  signal EQ_u16_u1_234_inst_ack_1 : boolean;
  signal type_cast_658_inst_req_1 : boolean;
  signal ULT_u16_u1_692_inst_req_0 : boolean;
  signal type_cast_658_inst_ack_1 : boolean;
  signal if_stmt_236_branch_req_0 : boolean;
  signal if_stmt_236_branch_ack_1 : boolean;
  signal if_stmt_236_branch_ack_0 : boolean;
  signal ADD_u16_u16_257_inst_req_0 : boolean;
  signal ADD_u16_u16_257_inst_ack_0 : boolean;
  signal ADD_u16_u16_257_inst_req_1 : boolean;
  signal ADD_u16_u16_257_inst_ack_1 : boolean;
  signal ADD_u16_u16_263_inst_req_0 : boolean;
  signal ADD_u16_u16_263_inst_ack_0 : boolean;
  signal ADD_u16_u16_263_inst_req_1 : boolean;
  signal ADD_u16_u16_263_inst_ack_1 : boolean;
  signal LOAD_ncol_ind_266_load_0_req_0 : boolean;
  signal LOAD_ncol_ind_266_load_0_ack_0 : boolean;
  signal LOAD_ncol_ind_266_load_0_req_1 : boolean;
  signal LOAD_ncol_ind_266_load_0_ack_1 : boolean;
  signal type_cast_271_inst_req_0 : boolean;
  signal type_cast_271_inst_ack_0 : boolean;
  signal type_cast_271_inst_req_1 : boolean;
  signal type_cast_271_inst_ack_1 : boolean;
  signal LOAD_nrows_274_load_0_req_0 : boolean;
  signal LOAD_nrows_274_load_0_ack_0 : boolean;
  signal LOAD_nrows_274_load_0_req_1 : boolean;
  signal LOAD_nrows_274_load_0_ack_1 : boolean;
  signal type_cast_278_inst_req_0 : boolean;
  signal type_cast_278_inst_ack_0 : boolean;
  signal type_cast_278_inst_req_1 : boolean;
  signal type_cast_278_inst_ack_1 : boolean;
  signal ADD_u32_u32_284_inst_req_0 : boolean;
  signal ADD_u32_u32_284_inst_ack_0 : boolean;
  signal ADD_u32_u32_284_inst_req_1 : boolean;
  signal ADD_u32_u32_284_inst_ack_1 : boolean;
  signal EQ_u32_u1_289_inst_req_0 : boolean;
  signal EQ_u32_u1_289_inst_ack_0 : boolean;
  signal EQ_u32_u1_289_inst_req_1 : boolean;
  signal EQ_u32_u1_289_inst_ack_1 : boolean;
  signal type_cast_293_inst_req_0 : boolean;
  signal type_cast_293_inst_ack_0 : boolean;
  signal type_cast_293_inst_req_1 : boolean;
  signal type_cast_293_inst_ack_1 : boolean;
  signal type_cast_297_inst_req_0 : boolean;
  signal type_cast_297_inst_ack_0 : boolean;
  signal type_cast_297_inst_req_1 : boolean;
  signal type_cast_297_inst_ack_1 : boolean;
  signal ADD_u64_u64_403_inst_req_1 : boolean;
  signal ADD_u64_u64_403_inst_ack_1 : boolean;
  signal if_stmt_680_branch_req_0 : boolean;
  signal ADD_u64_u64_408_inst_req_0 : boolean;
  signal ADD_u64_u64_408_inst_ack_0 : boolean;
  signal ADD_u64_u64_408_inst_req_1 : boolean;
  signal ADD_u64_u64_408_inst_ack_1 : boolean;
  signal ptr_deref_666_store_0_ack_1 : boolean;
  signal ptr_deref_666_store_0_req_1 : boolean;
  signal addr_of_413_final_reg_req_0 : boolean;
  signal addr_of_413_final_reg_ack_0 : boolean;
  signal addr_of_413_final_reg_req_1 : boolean;
  signal addr_of_413_final_reg_ack_1 : boolean;
  signal EQ_u16_u1_678_inst_ack_1 : boolean;
  signal EQ_u16_u1_678_inst_req_1 : boolean;
  signal ptr_deref_666_store_0_ack_0 : boolean;
  signal EQ_u16_u1_678_inst_ack_0 : boolean;
  signal EQ_u16_u1_678_inst_req_0 : boolean;
  signal ptr_deref_666_store_0_req_0 : boolean;
  signal ptr_deref_417_load_0_req_0 : boolean;
  signal ptr_deref_417_load_0_ack_0 : boolean;
  signal ptr_deref_417_load_0_req_1 : boolean;
  signal ptr_deref_417_load_0_ack_1 : boolean;
  signal type_cast_658_inst_ack_0 : boolean;
  signal ADD_u16_u16_423_inst_req_0 : boolean;
  signal ADD_u16_u16_423_inst_ack_0 : boolean;
  signal ADD_u16_u16_423_inst_req_1 : boolean;
  signal ADD_u16_u16_423_inst_ack_1 : boolean;
  signal type_cast_658_inst_req_0 : boolean;
  signal ADD_u16_u16_438_inst_req_0 : boolean;
  signal ADD_u16_u16_438_inst_ack_0 : boolean;
  signal ADD_u16_u16_438_inst_req_1 : boolean;
  signal ADD_u16_u16_438_inst_ack_1 : boolean;
  signal ADD_u16_u16_475_inst_req_0 : boolean;
  signal ADD_u16_u16_475_inst_ack_0 : boolean;
  signal ADD_u16_u16_475_inst_req_1 : boolean;
  signal ADD_u16_u16_475_inst_ack_1 : boolean;
  signal ADD_u16_u16_673_inst_ack_1 : boolean;
  signal type_cast_479_inst_req_0 : boolean;
  signal type_cast_479_inst_ack_0 : boolean;
  signal type_cast_479_inst_req_1 : boolean;
  signal type_cast_479_inst_ack_1 : boolean;
  signal ADD_u16_u16_673_inst_req_1 : boolean;
  signal addr_of_484_final_reg_req_0 : boolean;
  signal addr_of_484_final_reg_ack_0 : boolean;
  signal addr_of_484_final_reg_req_1 : boolean;
  signal addr_of_484_final_reg_ack_1 : boolean;
  signal ptr_deref_488_load_0_req_0 : boolean;
  signal ptr_deref_488_load_0_ack_0 : boolean;
  signal addr_of_663_final_reg_ack_1 : boolean;
  signal ptr_deref_488_load_0_req_1 : boolean;
  signal ptr_deref_488_load_0_ack_1 : boolean;
  signal addr_of_663_final_reg_req_1 : boolean;
  signal type_cast_492_inst_req_0 : boolean;
  signal type_cast_492_inst_ack_0 : boolean;
  signal type_cast_492_inst_req_1 : boolean;
  signal type_cast_492_inst_ack_1 : boolean;
  signal addr_of_663_final_reg_ack_0 : boolean;
  signal SLT_f64_u1_498_inst_req_0 : boolean;
  signal SLT_f64_u1_498_inst_ack_0 : boolean;
  signal SLT_f64_u1_498_inst_req_1 : boolean;
  signal SLT_f64_u1_498_inst_ack_1 : boolean;
  signal if_stmt_500_branch_req_0 : boolean;
  signal if_stmt_500_branch_ack_1 : boolean;
  signal if_stmt_500_branch_ack_0 : boolean;
  signal SUB_f32_f32_511_inst_req_0 : boolean;
  signal SUB_f32_f32_511_inst_ack_0 : boolean;
  signal SUB_f32_f32_511_inst_req_1 : boolean;
  signal SUB_f32_f32_511_inst_ack_1 : boolean;
  signal EQ_u16_u1_525_inst_req_0 : boolean;
  signal EQ_u16_u1_525_inst_ack_0 : boolean;
  signal EQ_u16_u1_525_inst_req_1 : boolean;
  signal EQ_u16_u1_525_inst_ack_1 : boolean;
  signal if_stmt_527_branch_req_0 : boolean;
  signal if_stmt_527_branch_ack_1 : boolean;
  signal if_stmt_527_branch_ack_0 : boolean;
  signal SLT_f64_u1_538_inst_req_0 : boolean;
  signal SLT_f64_u1_538_inst_ack_0 : boolean;
  signal SLT_f64_u1_538_inst_req_1 : boolean;
  signal SLT_f64_u1_538_inst_ack_1 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal type_cast_542_inst_req_1 : boolean;
  signal type_cast_542_inst_ack_1 : boolean;
  signal XOR_u8_u8_547_inst_req_0 : boolean;
  signal XOR_u8_u8_547_inst_ack_0 : boolean;
  signal XOR_u8_u8_547_inst_req_1 : boolean;
  signal XOR_u8_u8_547_inst_ack_1 : boolean;
  signal EQ_u8_u1_553_inst_req_0 : boolean;
  signal EQ_u8_u1_553_inst_ack_0 : boolean;
  signal EQ_u8_u1_553_inst_req_1 : boolean;
  signal EQ_u8_u1_553_inst_ack_1 : boolean;
  signal if_stmt_555_branch_req_0 : boolean;
  signal if_stmt_555_branch_ack_1 : boolean;
  signal if_stmt_555_branch_ack_0 : boolean;
  signal SLT_f32_u1_565_inst_req_0 : boolean;
  signal SLT_f32_u1_565_inst_ack_0 : boolean;
  signal SLT_f32_u1_565_inst_req_1 : boolean;
  signal SLT_f32_u1_565_inst_ack_1 : boolean;
  signal if_stmt_567_branch_req_0 : boolean;
  signal if_stmt_567_branch_ack_1 : boolean;
  signal if_stmt_567_branch_ack_0 : boolean;
  signal ADD_u16_u16_614_inst_req_0 : boolean;
  signal ADD_u16_u16_614_inst_ack_0 : boolean;
  signal ADD_u16_u16_614_inst_req_1 : boolean;
  signal ADD_u16_u16_614_inst_ack_1 : boolean;
  signal EQ_u16_u1_619_inst_req_0 : boolean;
  signal EQ_u16_u1_619_inst_ack_0 : boolean;
  signal EQ_u16_u1_619_inst_req_1 : boolean;
  signal EQ_u16_u1_619_inst_ack_1 : boolean;
  signal if_stmt_621_branch_req_0 : boolean;
  signal if_stmt_621_branch_ack_1 : boolean;
  signal if_stmt_621_branch_ack_0 : boolean;
  signal EQ_u8_u1_641_inst_req_0 : boolean;
  signal EQ_u8_u1_641_inst_ack_0 : boolean;
  signal EQ_u8_u1_641_inst_req_1 : boolean;
  signal EQ_u8_u1_641_inst_ack_1 : boolean;
  signal MUX_649_inst_req_0 : boolean;
  signal MUX_649_inst_ack_0 : boolean;
  signal MUX_649_inst_req_1 : boolean;
  signal MUX_649_inst_ack_1 : boolean;
  signal MUL_f32_f32_654_inst_req_0 : boolean;
  signal MUL_f32_f32_654_inst_ack_0 : boolean;
  signal MUL_f32_f32_654_inst_req_1 : boolean;
  signal MUL_f32_f32_654_inst_ack_1 : boolean;
  signal ULT_u16_u1_692_inst_req_1 : boolean;
  signal ULT_u16_u1_692_inst_ack_1 : boolean;
  signal if_stmt_694_branch_req_0 : boolean;
  signal if_stmt_694_branch_ack_1 : boolean;
  signal if_stmt_694_branch_ack_0 : boolean;
  signal phi_stmt_245_req_1 : boolean;
  signal type_cast_248_inst_req_0 : boolean;
  signal type_cast_248_inst_ack_0 : boolean;
  signal type_cast_248_inst_req_1 : boolean;
  signal type_cast_248_inst_ack_1 : boolean;
  signal phi_stmt_245_req_0 : boolean;
  signal phi_stmt_245_ack_0 : boolean;
  signal type_cast_378_inst_req_0 : boolean;
  signal type_cast_378_inst_ack_0 : boolean;
  signal type_cast_378_inst_req_1 : boolean;
  signal type_cast_378_inst_ack_1 : boolean;
  signal phi_stmt_375_req_0 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal phi_stmt_375_req_1 : boolean;
  signal phi_stmt_375_ack_0 : boolean;
  signal phi_stmt_427_req_0 : boolean;
  signal type_cast_433_inst_req_0 : boolean;
  signal type_cast_433_inst_ack_0 : boolean;
  signal type_cast_433_inst_req_1 : boolean;
  signal type_cast_433_inst_ack_1 : boolean;
  signal phi_stmt_427_req_1 : boolean;
  signal phi_stmt_427_ack_0 : boolean;
  signal type_cast_449_inst_req_0 : boolean;
  signal type_cast_449_inst_ack_0 : boolean;
  signal type_cast_449_inst_req_1 : boolean;
  signal type_cast_449_inst_ack_1 : boolean;
  signal phi_stmt_442_req_1 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal phi_stmt_450_req_1 : boolean;
  signal type_cast_463_inst_req_0 : boolean;
  signal type_cast_463_inst_ack_0 : boolean;
  signal type_cast_463_inst_req_1 : boolean;
  signal type_cast_463_inst_ack_1 : boolean;
  signal phi_stmt_457_req_1 : boolean;
  signal type_cast_470_inst_req_0 : boolean;
  signal type_cast_470_inst_ack_0 : boolean;
  signal type_cast_470_inst_req_1 : boolean;
  signal type_cast_470_inst_ack_1 : boolean;
  signal phi_stmt_464_req_1 : boolean;
  signal phi_stmt_442_req_0 : boolean;
  signal phi_stmt_450_req_0 : boolean;
  signal phi_stmt_457_req_0 : boolean;
  signal phi_stmt_464_req_0 : boolean;
  signal phi_stmt_442_ack_0 : boolean;
  signal phi_stmt_450_ack_0 : boolean;
  signal phi_stmt_457_ack_0 : boolean;
  signal phi_stmt_464_ack_0 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal phi_stmt_515_req_1 : boolean;
  signal type_cast_518_inst_req_0 : boolean;
  signal type_cast_518_inst_ack_0 : boolean;
  signal type_cast_518_inst_req_1 : boolean;
  signal type_cast_518_inst_ack_1 : boolean;
  signal phi_stmt_515_req_0 : boolean;
  signal phi_stmt_515_ack_0 : boolean;
  signal type_cast_579_inst_req_0 : boolean;
  signal type_cast_579_inst_ack_0 : boolean;
  signal type_cast_579_inst_req_1 : boolean;
  signal type_cast_579_inst_ack_1 : boolean;
  signal phi_stmt_576_req_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal phi_stmt_589_req_0 : boolean;
  signal type_cast_602_inst_req_0 : boolean;
  signal type_cast_602_inst_ack_0 : boolean;
  signal type_cast_602_inst_req_1 : boolean;
  signal type_cast_602_inst_ack_1 : boolean;
  signal phi_stmt_599_req_0 : boolean;
  signal phi_stmt_576_req_1 : boolean;
  signal type_cast_594_inst_req_0 : boolean;
  signal type_cast_594_inst_ack_0 : boolean;
  signal type_cast_594_inst_req_1 : boolean;
  signal type_cast_594_inst_ack_1 : boolean;
  signal phi_stmt_589_req_1 : boolean;
  signal type_cast_604_inst_req_0 : boolean;
  signal type_cast_604_inst_ack_0 : boolean;
  signal type_cast_604_inst_req_1 : boolean;
  signal type_cast_604_inst_ack_1 : boolean;
  signal phi_stmt_599_req_1 : boolean;
  signal phi_stmt_576_req_3 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal phi_stmt_589_req_3 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal phi_stmt_599_req_3 : boolean;
  signal phi_stmt_576_req_2 : boolean;
  signal type_cast_596_inst_req_0 : boolean;
  signal type_cast_596_inst_ack_0 : boolean;
  signal type_cast_596_inst_req_1 : boolean;
  signal type_cast_596_inst_ack_1 : boolean;
  signal phi_stmt_589_req_2 : boolean;
  signal type_cast_606_inst_req_0 : boolean;
  signal type_cast_606_inst_ack_0 : boolean;
  signal type_cast_606_inst_req_1 : boolean;
  signal type_cast_606_inst_ack_1 : boolean;
  signal phi_stmt_599_req_2 : boolean;
  signal phi_stmt_576_ack_0 : boolean;
  signal phi_stmt_589_ack_0 : boolean;
  signal phi_stmt_599_ack_0 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal phi_stmt_628_req_0 : boolean;
  signal type_cast_635_inst_req_0 : boolean;
  signal type_cast_635_inst_ack_0 : boolean;
  signal type_cast_635_inst_req_1 : boolean;
  signal type_cast_635_inst_ack_1 : boolean;
  signal phi_stmt_632_req_0 : boolean;
  signal phi_stmt_628_ack_0 : boolean;
  signal phi_stmt_632_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "checkNodeComputeEngine_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  checkNodeComputeEngine_CP_1062_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "checkNodeComputeEngine_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= checkNodeComputeEngine_CP_1062_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= checkNodeComputeEngine_CP_1062_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= checkNodeComputeEngine_CP_1062_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  checkNodeComputeEngine_CP_1062: Block -- control-path 
    signal checkNodeComputeEngine_CP_1062_elements: BooleanArray(442 downto 0);
    -- 
  begin -- 
    checkNodeComputeEngine_CP_1062_elements(0) <= checkNodeComputeEngine_CP_1062_start;
    checkNodeComputeEngine_CP_1062_symbol <= checkNodeComputeEngine_CP_1062_elements(442);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_226/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	37 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_226/branch_block_stmt_226__entry__
      -- CP-element group 1: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(1) <= checkNodeComputeEngine_CP_1062_elements(0);
    -- CP-element group 2:  branch  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	41 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	42 
    -- CP-element group 2: 	43 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235__exit__
      -- CP-element group 2: 	 branch_block_stmt_226/if_stmt_236__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(2) <= checkNodeComputeEngine_CP_1062_elements(41);
    -- CP-element group 3:  merge  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	270 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	271 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_226/merge_stmt_242__exit__
      -- CP-element group 3: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11
      -- 
    checkNodeComputeEngine_CP_1062_elements(3) <= checkNodeComputeEngine_CP_1062_elements(270);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	280 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	51 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_226/merge_stmt_244__exit__
      -- CP-element group 4: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(4) <= checkNodeComputeEngine_CP_1062_elements(280);
    -- CP-element group 5:  branch  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	78 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	79 
    -- CP-element group 5: 	80 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309__exit__
      -- CP-element group 5: 	 branch_block_stmt_226/if_stmt_310__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(5) <= checkNodeComputeEngine_CP_1062_elements(78);
    -- CP-element group 6:  merge  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	283 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	88 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_226/merge_stmt_316__exit__
      -- CP-element group 6: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(6) <= checkNodeComputeEngine_CP_1062_elements(283);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	104 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	291 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350__exit__
      -- CP-element group 7: 	 branch_block_stmt_226/bb_4_bb_5
      -- 
    checkNodeComputeEngine_CP_1062_elements(7) <= checkNodeComputeEngine_CP_1062_elements(104);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	286 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	105 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_226/merge_stmt_352__exit__
      -- CP-element group 8: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(8) <= checkNodeComputeEngine_CP_1062_elements(286);
    -- CP-element group 9:  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	115 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	287 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372__exit__
      -- CP-element group 9: 	 branch_block_stmt_226/bb_3_bb_5
      -- 
    checkNodeComputeEngine_CP_1062_elements(9) <= checkNodeComputeEngine_CP_1062_elements(115);
    -- CP-element group 10:  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	297 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	116 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_226/merge_stmt_374__exit__
      -- CP-element group 10: 	 branch_block_stmt_226/assign_stmt_387__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(10) <= checkNodeComputeEngine_CP_1062_elements(297);
    -- CP-element group 11:  branch  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	118 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	120 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_226/assign_stmt_387__exit__
      -- CP-element group 11: 	 branch_block_stmt_226/if_stmt_388__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(11) <= checkNodeComputeEngine_CP_1062_elements(118);
    -- CP-element group 12:  merge  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	300 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	128 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_226/merge_stmt_394__exit__
      -- CP-element group 12: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(12) <= checkNodeComputeEngine_CP_1062_elements(300);
    -- CP-element group 13:  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	141 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	301 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424__exit__
      -- CP-element group 13: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph
      -- 
    checkNodeComputeEngine_CP_1062_elements(13) <= checkNodeComputeEngine_CP_1062_elements(141);
    -- CP-element group 14:  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	310 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	142 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_226/merge_stmt_426__exit__
      -- CP-element group 14: 	 branch_block_stmt_226/assign_stmt_439__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(14) <= checkNodeComputeEngine_CP_1062_elements(310);
    -- CP-element group 15:  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	144 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	325 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_226/assign_stmt_439__exit__
      -- CP-element group 15: 	 branch_block_stmt_226/bbx_xnph_bb_8
      -- 
    checkNodeComputeEngine_CP_1062_elements(15) <= checkNodeComputeEngine_CP_1062_elements(144);
    -- CP-element group 16:  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	341 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	145 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_226/merge_stmt_441__exit__
      -- CP-element group 16: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(16) <= checkNodeComputeEngine_CP_1062_elements(341);
    -- CP-element group 17:  branch  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	158 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	159 
    -- CP-element group 17: 	160 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499__exit__
      -- CP-element group 17: 	 branch_block_stmt_226/if_stmt_500__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(17) <= checkNodeComputeEngine_CP_1062_elements(158);
    -- CP-element group 18:  merge  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	344 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	168 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_226/merge_stmt_506__exit__
      -- CP-element group 18: 	 branch_block_stmt_226/assign_stmt_512__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(18) <= checkNodeComputeEngine_CP_1062_elements(344);
    -- CP-element group 19:  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	170 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	349 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_226/assign_stmt_512__exit__
      -- CP-element group 19: 	 branch_block_stmt_226/bb_9_bb_10
      -- 
    checkNodeComputeEngine_CP_1062_elements(19) <= checkNodeComputeEngine_CP_1062_elements(170);
    -- CP-element group 20:  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	355 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	171 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_226/merge_stmt_514__exit__
      -- CP-element group 20: 	 branch_block_stmt_226/assign_stmt_526__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(20) <= checkNodeComputeEngine_CP_1062_elements(355);
    -- CP-element group 21:  branch  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	173 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	174 
    -- CP-element group 21: 	175 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_226/assign_stmt_526__exit__
      -- CP-element group 21: 	 branch_block_stmt_226/if_stmt_527__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(21) <= checkNodeComputeEngine_CP_1062_elements(173);
    -- CP-element group 22:  merge  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	358 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	183 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_226/merge_stmt_533__exit__
      -- CP-element group 22: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(22) <= checkNodeComputeEngine_CP_1062_elements(358);
    -- CP-element group 23:  branch  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	192 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	193 
    -- CP-element group 23: 	194 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554__exit__
      -- CP-element group 23: 	 branch_block_stmt_226/if_stmt_555__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(23) <= checkNodeComputeEngine_CP_1062_elements(192);
    -- CP-element group 24:  merge  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	361 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	202 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_226/merge_stmt_561__exit__
      -- CP-element group 24: 	 branch_block_stmt_226/assign_stmt_566__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(24) <= checkNodeComputeEngine_CP_1062_elements(361);
    -- CP-element group 25:  branch  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	204 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	205 
    -- CP-element group 25: 	206 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_226/assign_stmt_566__exit__
      -- CP-element group 25: 	 branch_block_stmt_226/if_stmt_567__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(25) <= checkNodeComputeEngine_CP_1062_elements(204);
    -- CP-element group 26:  merge  place  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	364 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	396 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_226/merge_stmt_573__exit__
      -- CP-element group 26: 	 branch_block_stmt_226/bb_13_bb_14
      -- 
    checkNodeComputeEngine_CP_1062_elements(26) <= checkNodeComputeEngine_CP_1062_elements(364);
    -- CP-element group 27:  place  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	411 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	214 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_226/merge_stmt_575__exit__
      -- CP-element group 27: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(27) <= checkNodeComputeEngine_CP_1062_elements(411);
    -- CP-element group 28:  branch  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	218 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	219 
    -- CP-element group 28: 	220 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620__exit__
      -- CP-element group 28: 	 branch_block_stmt_226/if_stmt_621__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(28) <= checkNodeComputeEngine_CP_1062_elements(218);
    -- CP-element group 29:  merge  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	424 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	228 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_226/merge_stmt_627__exit__
      -- CP-element group 29: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(29) <= checkNodeComputeEngine_CP_1062_elements(424);
    -- CP-element group 30:  branch  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	246 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	247 
    -- CP-element group 30: 	248 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679__exit__
      -- CP-element group 30: 	 branch_block_stmt_226/if_stmt_680__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(30) <= checkNodeComputeEngine_CP_1062_elements(246);
    -- CP-element group 31:  merge  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	427 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	429 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_226/merge_stmt_686__exit__
      -- CP-element group 31: 	 branch_block_stmt_226/xx_x_crit_edge9x_xloopexit_xx_x_crit_edge9
      -- 
    checkNodeComputeEngine_CP_1062_elements(31) <= checkNodeComputeEngine_CP_1062_elements(427);
    -- CP-element group 32:  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	431 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	256 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_226/merge_stmt_688__exit__
      -- CP-element group 32: 	 branch_block_stmt_226/assign_stmt_693__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(32) <= checkNodeComputeEngine_CP_1062_elements(431);
    -- CP-element group 33:  branch  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	258 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	259 
    -- CP-element group 33: 	260 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_226/assign_stmt_693__exit__
      -- CP-element group 33: 	 branch_block_stmt_226/if_stmt_694__entry__
      -- 
    checkNodeComputeEngine_CP_1062_elements(33) <= checkNodeComputeEngine_CP_1062_elements(258);
    -- CP-element group 34:  merge  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	434 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	436 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_226/merge_stmt_700__exit__
      -- CP-element group 34: 	 branch_block_stmt_226/xx_x_crit_edge12x_xloopexit_xx_x_crit_edge12
      -- 
    checkNodeComputeEngine_CP_1062_elements(34) <= checkNodeComputeEngine_CP_1062_elements(434);
    -- CP-element group 35:  place  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	438 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	439 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_226/merge_stmt_702__exit__
      -- CP-element group 35: 	 branch_block_stmt_226/return__
      -- 
    checkNodeComputeEngine_CP_1062_elements(35) <= checkNodeComputeEngine_CP_1062_elements(438);
    -- CP-element group 36:  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	441 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	442 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_226/branch_block_stmt_226__exit__
      -- CP-element group 36: 	 branch_block_stmt_226/merge_stmt_704__exit__
      -- 
    checkNodeComputeEngine_CP_1062_elements(36) <= checkNodeComputeEngine_CP_1062_elements(441);
    -- CP-element group 37:  fork  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	1 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	41 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_update_start_
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/word_0/rr
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_update_start_
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Update/cr
      -- 
    cr_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(37), ack => LOAD_nrows_228_load_0_req_1); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(37), ack => LOAD_nrows_228_load_0_req_0); -- 
    cr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(37), ack => EQ_u16_u1_234_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(37) <= checkNodeComputeEngine_CP_1062_elements(1);
    -- CP-element group 38:  transition  input  no-bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Sample/word_access_start/word_0/ra
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_228_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  no-bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (12) 
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/LOAD_nrows_228_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/LOAD_nrows_228_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/LOAD_nrows_228_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/LOAD_nrows_228_Update/LOAD_nrows_228_Merge/merge_ack
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Sample/rr
      -- 
    ca_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_228_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(39)); -- 
    rr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(39), ack => EQ_u16_u1_234_inst_req_0); -- 
    -- CP-element group 40:  transition  input  no-bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Sample/ra
      -- 
    ra_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_234_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(40)); -- 
    -- CP-element group 41:  transition  input  no-bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	37 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	2 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/$exit
      -- CP-element group 41: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_226/assign_stmt_229_to_assign_stmt_235/EQ_u16_u1_234_Update/ca
      -- 
    ca_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_234_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(41)); -- 
    -- CP-element group 42:  transition  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	2 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_226/if_stmt_236_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(42) <= checkNodeComputeEngine_CP_1062_elements(2);
    -- CP-element group 43:  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	2 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_226/if_stmt_236_eval_test/$entry
      -- CP-element group 43: 	 branch_block_stmt_226/if_stmt_236_eval_test/$exit
      -- CP-element group 43: 	 branch_block_stmt_226/if_stmt_236_eval_test/branch_req
      -- 
    branch_req_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(43), ack => if_stmt_236_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(43) <= checkNodeComputeEngine_CP_1062_elements(2);
    -- CP-element group 44:  branch  place  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_226/R_iNsTr_1_237_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(44) <= checkNodeComputeEngine_CP_1062_elements(43);
    -- CP-element group 45:  transition  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_226/if_stmt_236_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(45) <= checkNodeComputeEngine_CP_1062_elements(44);
    -- CP-element group 46:  transition  input  no-bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_226/if_stmt_236_if_link/$exit
      -- CP-element group 46: 	 branch_block_stmt_226/if_stmt_236_if_link/if_choice_transition
      -- 
    if_choice_transition_1222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_236_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(46)); -- 
    -- CP-element group 47:  transition  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_226/if_stmt_236_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(47) <= checkNodeComputeEngine_CP_1062_elements(44);
    -- CP-element group 48:  transition  input  no-bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_226/if_stmt_236_else_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_226/if_stmt_236_else_link/else_choice_transition
      -- 
    else_choice_transition_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_236_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(48)); -- 
    -- CP-element group 49:  place  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	435 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_226/bb_0_xx_x_crit_edge12
      -- 
    checkNodeComputeEngine_CP_1062_elements(49) <= checkNodeComputeEngine_CP_1062_elements(46);
    -- CP-element group 50:  place  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	268 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_226/bb_0_bbx_xnph11x_xpreheader
      -- 
    checkNodeComputeEngine_CP_1062_elements(50) <= checkNodeComputeEngine_CP_1062_elements(48);
    -- CP-element group 51:  fork  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	4 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	55 
    -- CP-element group 51: 	56 
    -- CP-element group 51: 	57 
    -- CP-element group 51: 	58 
    -- CP-element group 51: 	59 
    -- CP-element group 51: 	60 
    -- CP-element group 51: 	61 
    -- CP-element group 51: 	63 
    -- CP-element group 51: 	65 
    -- CP-element group 51: 	68 
    -- CP-element group 51: 	70 
    -- CP-element group 51: 	71 
    -- CP-element group 51: 	72 
    -- CP-element group 51: 	74 
    -- CP-element group 51: 	77 
    -- CP-element group 51:  members (67) 
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/word_0/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/word_0/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/word_0/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/word_0/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_update_start_
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Update/cr
      -- 
    rr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u16_u16_257_inst_req_0); -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u16_u16_257_inst_req_1); -- 
    rr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u16_u16_263_inst_req_0); -- 
    cr_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u16_u16_263_inst_req_1); -- 
    cr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => LOAD_ncol_ind_266_load_0_req_1); -- 
    rr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => LOAD_ncol_ind_266_load_0_req_0); -- 
    rr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_271_inst_req_0); -- 
    cr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_271_inst_req_1); -- 
    cr_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => LOAD_nrows_274_load_0_req_1); -- 
    rr_1322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => LOAD_nrows_274_load_0_req_0); -- 
    cr_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_278_inst_req_1); -- 
    cr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u32_u32_284_inst_req_1); -- 
    cr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => EQ_u32_u1_289_inst_req_1); -- 
    cr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_293_inst_req_1); -- 
    rr_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_297_inst_req_0); -- 
    cr_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => type_cast_297_inst_req_1); -- 
    cr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u64_u64_303_inst_req_1); -- 
    cr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(51), ack => ADD_u64_u64_308_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(51) <= checkNodeComputeEngine_CP_1062_elements(4);
    -- CP-element group 52:  transition  input  no-bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Sample/ra
      -- 
    ra_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_257_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(52)); -- 
    -- CP-element group 53:  transition  input  no-bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_257_Update/ca
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_257_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(53)); -- 
    -- CP-element group 54:  transition  input  no-bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Sample/ra
      -- 
    ra_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_263_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(54)); -- 
    -- CP-element group 55:  transition  input  no-bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	51 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	78 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u16_u16_263_Update/ca
      -- 
    ca_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_263_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(55)); -- 
    -- CP-element group 56:  transition  input  no-bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	51 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Sample/word_access_start/word_0/ra
      -- 
    ra_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_266_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  no-bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	69 
    -- CP-element group 57:  members (12) 
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/LOAD_ncol_ind_266_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/LOAD_ncol_ind_266_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/LOAD_ncol_ind_266_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_ncol_ind_266_Update/LOAD_ncol_ind_266_Merge/merge_ack
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Sample/rr
      -- 
    ca_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_266_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(57)); -- 
    rr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(57), ack => type_cast_293_inst_req_0); -- 
    -- CP-element group 58:  transition  input  no-bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Sample/ra
      -- 
    ra_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_271_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(58)); -- 
    -- CP-element group 59:  transition  input  no-bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	66 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_271_Update/ca
      -- 
    ca_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_271_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(59)); -- 
    -- CP-element group 60:  transition  input  no-bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	51 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/$exit
      -- CP-element group 60: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Sample/word_access_start/word_0/ra
      -- 
    ra_1323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_274_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  no-bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	51 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/$exit
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/word_0/$exit
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/word_access_complete/word_0/ca
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/LOAD_nrows_274_Merge/$entry
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/LOAD_nrows_274_Merge/$exit
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/LOAD_nrows_274_Merge/merge_req
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/LOAD_nrows_274_Update/LOAD_nrows_274_Merge/merge_ack
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Sample/rr
      -- 
    ca_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_274_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(61)); -- 
    rr_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(61), ack => type_cast_278_inst_req_0); -- 
    -- CP-element group 62:  transition  input  no-bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Sample/ra
      -- 
    ra_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_278_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  no-bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	51 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_278_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Sample/rr
      -- 
    ca_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_278_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(63)); -- 
    rr_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(63), ack => ADD_u32_u32_284_inst_req_0); -- 
    -- CP-element group 64:  transition  input  no-bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Sample/ra
      -- 
    ra_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_284_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(64)); -- 
    -- CP-element group 65:  transition  input  no-bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	51 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u32_u32_284_Update/ca
      -- 
    ca_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_284_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	59 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Sample/rr
      -- 
    rr_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(66), ack => EQ_u32_u1_289_inst_req_0); -- 
    checkNodeComputeEngine_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 42) := "checkNodeComputeEngine_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(59) & checkNodeComputeEngine_CP_1062_elements(65);
      gj_checkNodeComputeEngine_cp_element_group_66 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  no-bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Sample/ra
      -- 
    ra_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_289_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(67)); -- 
    -- CP-element group 68:  transition  input  no-bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	51 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	78 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/EQ_u32_u1_289_Update/ca
      -- 
    ca_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_289_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(68)); -- 
    -- CP-element group 69:  transition  input  no-bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	57 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Sample/ra
      -- 
    ra_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_293_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(69)); -- 
    -- CP-element group 70:  transition  input  no-bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	51 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_293_Update/ca
      -- 
    ca_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_293_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(70)); -- 
    -- CP-element group 71:  transition  input  no-bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	51 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Sample/ra
      -- 
    ra_1404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  no-bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	51 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/type_cast_297_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_sample_start_
      -- 
    ca_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(72)); -- 
    rr_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(72), ack => ADD_u64_u64_303_inst_req_0); -- 
    -- CP-element group 73:  transition  input  no-bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_sample_completed_
      -- 
    ra_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_303_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(73)); -- 
    -- CP-element group 74:  transition  input  no-bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	51 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_303_update_completed_
      -- 
    ca_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_303_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Sample/rr
      -- 
    rr_1431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(75), ack => ADD_u64_u64_308_inst_req_0); -- 
    checkNodeComputeEngine_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 42) := "checkNodeComputeEngine_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(70) & checkNodeComputeEngine_CP_1062_elements(74);
      gj_checkNodeComputeEngine_cp_element_group_75 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  no-bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Sample/ra
      -- 
    ra_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_308_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(76)); -- 
    -- CP-element group 77:  transition  input  no-bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	51 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/ADD_u64_u64_308_Update/ca
      -- 
    ca_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_308_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: 	55 
    -- CP-element group 78: 	68 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	5 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_226/assign_stmt_258_to_assign_stmt_309/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 42) := "checkNodeComputeEngine_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(53) & checkNodeComputeEngine_CP_1062_elements(55) & checkNodeComputeEngine_CP_1062_elements(68) & checkNodeComputeEngine_CP_1062_elements(77);
      gj_checkNodeComputeEngine_cp_element_group_78 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	5 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_226/if_stmt_310_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(79) <= checkNodeComputeEngine_CP_1062_elements(5);
    -- CP-element group 80:  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	5 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_226/if_stmt_310_eval_test/$entry
      -- CP-element group 80: 	 branch_block_stmt_226/if_stmt_310_eval_test/$exit
      -- CP-element group 80: 	 branch_block_stmt_226/if_stmt_310_eval_test/branch_req
      -- 
    branch_req_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(80), ack => if_stmt_310_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(80) <= checkNodeComputeEngine_CP_1062_elements(5);
    -- CP-element group 81:  branch  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	84 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_226/R_iNsTr_13_311_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(81) <= checkNodeComputeEngine_CP_1062_elements(80);
    -- CP-element group 82:  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_226/if_stmt_310_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(82) <= checkNodeComputeEngine_CP_1062_elements(81);
    -- CP-element group 83:  transition  input  no-bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_226/if_stmt_310_if_link/$exit
      -- CP-element group 83: 	 branch_block_stmt_226/if_stmt_310_if_link/if_choice_transition
      -- 
    if_choice_transition_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_310_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(83)); -- 
    -- CP-element group 84:  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	81 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_226/if_stmt_310_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(84) <= checkNodeComputeEngine_CP_1062_elements(81);
    -- CP-element group 85:  transition  input  no-bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_226/if_stmt_310_else_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_226/if_stmt_310_else_link/else_choice_transition
      -- 
    else_choice_transition_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_310_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(85)); -- 
    -- CP-element group 86:  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	284 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_226/bbx_xnph11_bb_3
      -- 
    checkNodeComputeEngine_CP_1062_elements(86) <= checkNodeComputeEngine_CP_1062_elements(83);
    -- CP-element group 87:  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	281 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_226/bbx_xnph11_bb_4
      -- 
    checkNodeComputeEngine_CP_1062_elements(87) <= checkNodeComputeEngine_CP_1062_elements(85);
    -- CP-element group 88:  fork  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	6 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	90 
    -- CP-element group 88: 	92 
    -- CP-element group 88: 	93 
    -- CP-element group 88: 	94 
    -- CP-element group 88: 	96 
    -- CP-element group 88: 	98 
    -- CP-element group 88: 	100 
    -- CP-element group 88: 	103 
    -- CP-element group 88:  members (53) 
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_scale_0/scale_rename_req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_scaled_0
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_resize_0/index_resize_req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_resize_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_request/req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_resize_0/index_resize_ack
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_resize_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_resized_0
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_scale_0/scale_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_final_index_sum_regn/$exit
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_computed_0
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_final_index_sum_regn/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_final_index_sum_regn/req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_complete/req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_scale_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_final_index_sum_regn/ack
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_complete/req
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_330_index_scale_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_update_start_
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_update_start_
      -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => ADD_u64_u64_321_inst_req_0); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => ADD_u64_u64_321_inst_req_1); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => ADD_u64_u64_326_inst_req_1); -- 
    req_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => addr_of_331_final_reg_req_1); -- 
    req_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => addr_of_331_final_reg_req_0); -- 
    req_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => addr_of_336_final_reg_req_1); -- 
    cr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => ptr_deref_340_load_0_req_1); -- 
    cr_1659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => ptr_deref_344_load_0_req_1); -- 
    cr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(88), ack => SUB_u16_u16_349_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(88) <= checkNodeComputeEngine_CP_1062_elements(6);
    -- CP-element group 89:  transition  input  no-bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Sample/ra
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_321_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  no-bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_321_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_sample_start_
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_321_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(90)); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(90), ack => ADD_u64_u64_326_inst_req_0); -- 
    -- CP-element group 91:  transition  input  no-bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Sample/$exit
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_326_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  no-bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	88 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (27) 
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_computed_0
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_scaled_0
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_resize_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_scale_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_scale_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_base_plus_offset/$exit
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_scale_0/scale_rename_req
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_scale_0/scale_rename_ack
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_final_index_sum_regn/$entry
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_resize_0/index_resize_req
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_resize_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_final_index_sum_regn/$exit
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_resize_0/index_resize_ack
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_final_index_sum_regn/req
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_final_index_sum_regn/ack
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_base_plus_offset/$entry
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_base_plus_offset/sum_rename_req
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_base_plus_offset/sum_rename_ack
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_request/$entry
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_request/req
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ADD_u64_u64_326_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_index_resized_0
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_offset_calculated
      -- CP-element group 92: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/array_obj_ref_335_root_address_calculated
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_326_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(92)); -- 
    req_1559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(92), ack => addr_of_336_final_reg_req_0); -- 
    -- CP-element group 93:  transition  input  no-bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	88 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	104 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_request/$exit
      -- CP-element group 93: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_request/ack
      -- CP-element group 93: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_sample_completed_
      -- 
    ack_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_331_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(93)); -- 
    -- CP-element group 94:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	88 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	97 
    -- CP-element group 94:  members (24) 
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_addr_resize/$exit
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_word_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_root_address_calculated
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_address_resized
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_addr_resize/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_addr_resize/base_resize_req
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_addr_resize/base_resize_ack
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_plus_offset/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_plus_offset/$exit
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_plus_offset/sum_rename_req
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_base_plus_offset/sum_rename_ack
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_word_addrgen/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_word_addrgen/$exit
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_word_addrgen/root_register_req
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_word_addrgen/root_register_ack
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_331_complete/ack
      -- CP-element group 94: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_sample_start_
      -- 
    ack_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_331_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(94)); -- 
    rr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(94), ack => ptr_deref_340_load_0_req_0); -- 
    -- CP-element group 95:  transition  input  no-bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	104 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_request/$exit
      -- CP-element group 95: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_request/ack
      -- CP-element group 95: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_sample_completed_
      -- 
    ack_1560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_336_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	88 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (24) 
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_word_addrgen/root_register_req
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_word_addrgen/root_register_ack
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_word_addrgen/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/word_0/rr
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_word_addrgen/$exit
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_word_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_root_address_calculated
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_address_resized
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_addr_resize/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_addr_resize/$exit
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_addr_resize/base_resize_req
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_addr_resize/base_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_plus_offset/$entry
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_plus_offset/$exit
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_plus_offset/sum_rename_req
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_base_plus_offset/sum_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_complete/ack
      -- CP-element group 96: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/addr_of_336_update_completed_
      -- 
    ack_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_336_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(96)); -- 
    rr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(96), ack => ptr_deref_344_load_0_req_0); -- 
    -- CP-element group 97:  transition  input  no-bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	94 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Sample/word_access_start/word_0/ra
      -- CP-element group 97: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_sample_completed_
      -- 
    ra_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_340_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(97)); -- 
    -- CP-element group 98:  transition  input  no-bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	101 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/ptr_deref_340_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/ptr_deref_340_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/ptr_deref_340_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_340_Update/ptr_deref_340_Merge/merge_ack
      -- 
    ca_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_340_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(98)); -- 
    -- CP-element group 99:  transition  input  no-bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_sample_completed_
      -- 
    ra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_344_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(99)); -- 
    -- CP-element group 100:  transition  input  no-bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	88 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/ptr_deref_344_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/ptr_deref_344_Merge/$exit
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/ptr_deref_344_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_Update/ptr_deref_344_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/ptr_deref_344_update_completed_
      -- 
    ca_1660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_344_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	98 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Sample/rr
      -- 
    rr_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(101), ack => SUB_u16_u16_349_inst_req_0); -- 
    checkNodeComputeEngine_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(98) & checkNodeComputeEngine_CP_1062_elements(100);
      gj_checkNodeComputeEngine_cp_element_group_101 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  no-bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Sample/$exit
      -- 
    ra_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_349_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(102)); -- 
    -- CP-element group 103:  transition  input  no-bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	88 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/SUB_u16_u16_349_update_completed_
      -- 
    ca_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_349_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(103)); -- 
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	93 
    -- CP-element group 104: 	95 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	7 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_226/assign_stmt_322_to_assign_stmt_350/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(93) & checkNodeComputeEngine_CP_1062_elements(95) & checkNodeComputeEngine_CP_1062_elements(103);
      gj_checkNodeComputeEngine_cp_element_group_104 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	109 
    -- CP-element group 105: 	110 
    -- CP-element group 105: 	111 
    -- CP-element group 105: 	114 
    -- CP-element group 105:  members (42) 
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_update_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_resize_0/index_resize_ack
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_update_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/word_0/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_scale_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_final_index_sum_regn/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/word_0/cr
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_update_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_request/req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_update_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_scale_0/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_complete/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_final_index_sum_regn/$exit
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_final_index_sum_regn/req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_final_index_sum_regn/ack
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_base_plus_offset/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_complete/req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_scale_0/scale_rename_req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_base_plus_offset/$exit
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_base_plus_offset/sum_rename_req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_base_plus_offset/sum_rename_ack
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_scale_0/scale_rename_ack
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_request/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_resize_0/index_resize_req
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_resize_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_resize_0/$entry
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_computed_0
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_scaled_0
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_index_resized_0
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_offset_calculated
      -- CP-element group 105: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/array_obj_ref_355_root_address_calculated
      -- 
    req_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => addr_of_356_final_reg_req_1); -- 
    req_1715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => addr_of_356_final_reg_req_0); -- 
    cr_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => ptr_deref_360_load_0_req_1); -- 
    rr_1779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => ADD_u16_u16_366_inst_req_0); -- 
    cr_1784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => ADD_u16_u16_366_inst_req_1); -- 
    cr_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(105), ack => SUB_u16_u16_371_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(105) <= checkNodeComputeEngine_CP_1062_elements(8);
    -- CP-element group 106:  transition  input  no-bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	115 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_request/ack
      -- CP-element group 106: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_request/$exit
      -- 
    ack_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_356_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (24) 
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_plus_offset/sum_rename_req
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/$entry
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_root_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_plus_offset/$entry
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_addr_resize/$entry
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_word_addrgen/root_register_req
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/word_0/$entry
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_addr_resize/base_resize_ack
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_word_addrgen/root_register_ack
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/word_0/rr
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_plus_offset/$exit
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_addr_resize/$exit
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_word_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_address_resized
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_addr_resize/base_resize_req
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_complete/ack
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/addr_of_356_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_base_plus_offset/sum_rename_ack
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_word_addrgen/$exit
      -- CP-element group 107: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_word_addrgen/$entry
      -- 
    ack_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_356_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(107)); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(107), ack => ptr_deref_360_load_0_req_0); -- 
    -- CP-element group 108:  transition  input  no-bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/$exit
      -- CP-element group 108: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Sample/word_access_start/word_0/ra
      -- 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_360_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(108)); -- 
    -- CP-element group 109:  transition  input  no-bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	105 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/$exit
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/word_access_complete/word_0/ca
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/ptr_deref_360_Merge/$entry
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/ptr_deref_360_Merge/$exit
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/ptr_deref_360_Merge/merge_req
      -- CP-element group 109: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ptr_deref_360_Update/ptr_deref_360_Merge/merge_ack
      -- 
    ca_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_360_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(109)); -- 
    -- CP-element group 110:  transition  input  no-bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Sample/$exit
      -- 
    ra_1780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_366_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(110)); -- 
    -- CP-element group 111:  transition  input  no-bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	105 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/ADD_u16_u16_366_update_completed_
      -- 
    ca_1785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_366_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Sample/rr
      -- 
    rr_1793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(112), ack => SUB_u16_u16_371_inst_req_0); -- 
    checkNodeComputeEngine_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(109) & checkNodeComputeEngine_CP_1062_elements(111);
      gj_checkNodeComputeEngine_cp_element_group_112 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  no-bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Sample/ra
      -- 
    ra_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_371_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(113)); -- 
    -- CP-element group 114:  transition  input  no-bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	105 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/SUB_u16_u16_371_Update/ca
      -- 
    ca_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_371_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(114)); -- 
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	106 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	9 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_226/assign_stmt_357_to_assign_stmt_372/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(106) & checkNodeComputeEngine_CP_1062_elements(114);
      gj_checkNodeComputeEngine_cp_element_group_115 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	10 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (7) 
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_update_start_
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_226/assign_stmt_387/$entry
      -- 
    rr_1810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(116), ack => EQ_u16_u1_386_inst_req_0); -- 
    cr_1815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(116), ack => EQ_u16_u1_386_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(116) <= checkNodeComputeEngine_CP_1062_elements(10);
    -- CP-element group 117:  transition  input  no-bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Sample/$exit
      -- 
    ra_1811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_386_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(117)); -- 
    -- CP-element group 118:  transition  input  no-bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_226/assign_stmt_387/$exit
      -- CP-element group 118: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_226/assign_stmt_387/EQ_u16_u1_386_Update/ca
      -- 
    ca_1816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_386_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(118)); -- 
    -- CP-element group 119:  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	11 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_226/if_stmt_388_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(119) <= checkNodeComputeEngine_CP_1062_elements(11);
    -- CP-element group 120:  transition  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_226/if_stmt_388_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_226/if_stmt_388_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_226/if_stmt_388_eval_test/branch_req
      -- 
    branch_req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(120), ack => if_stmt_388_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(120) <= checkNodeComputeEngine_CP_1062_elements(11);
    -- CP-element group 121:  branch  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_226/R_iNsTr_31_389_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(121) <= checkNodeComputeEngine_CP_1062_elements(120);
    -- CP-element group 122:  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_226/if_stmt_388_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(122) <= checkNodeComputeEngine_CP_1062_elements(121);
    -- CP-element group 123:  transition  input  no-bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_226/if_stmt_388_if_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_226/if_stmt_388_if_link/if_choice_transition
      -- 
    if_choice_transition_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_388_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(123)); -- 
    -- CP-element group 124:  transition  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_226/if_stmt_388_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(124) <= checkNodeComputeEngine_CP_1062_elements(121);
    -- CP-element group 125:  transition  input  no-bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_226/if_stmt_388_else_link/else_choice_transition
      -- CP-element group 125: 	 branch_block_stmt_226/if_stmt_388_else_link/$exit
      -- 
    else_choice_transition_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_388_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(125)); -- 
    -- CP-element group 126:  place  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	428 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_226/bb_5_xx_x_crit_edge9
      -- 
    checkNodeComputeEngine_CP_1062_elements(126) <= checkNodeComputeEngine_CP_1062_elements(123);
    -- CP-element group 127:  place  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	298 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_226/bb_5_bbx_xnph8
      -- 
    checkNodeComputeEngine_CP_1062_elements(127) <= checkNodeComputeEngine_CP_1062_elements(125);
    -- CP-element group 128:  fork  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	12 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	130 
    -- CP-element group 128: 	132 
    -- CP-element group 128: 	134 
    -- CP-element group 128: 	136 
    -- CP-element group 128: 	138 
    -- CP-element group 128: 	140 
    -- CP-element group 128:  members (24) 
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Update/cr
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Update/cr
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Update/cr
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_complete/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_complete/req
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/word_0/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/word_0/cr
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_update_start_
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Update/cr
      -- 
    rr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => type_cast_397_inst_req_0); -- 
    cr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => type_cast_397_inst_req_1); -- 
    cr_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => ADD_u64_u64_403_inst_req_1); -- 
    cr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => ADD_u64_u64_408_inst_req_1); -- 
    req_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => addr_of_413_final_reg_req_1); -- 
    cr_1963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => ptr_deref_417_load_0_req_1); -- 
    cr_1982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(128), ack => ADD_u16_u16_423_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(128) <= checkNodeComputeEngine_CP_1062_elements(12);
    -- CP-element group 129:  transition  input  no-bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_sample_completed_
      -- 
    ra_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  no-bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/type_cast_397_update_completed_
      -- 
    ca_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(130)); -- 
    rr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(130), ack => ADD_u64_u64_403_inst_req_0); -- 
    -- CP-element group 131:  transition  input  no-bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_sample_completed_
      -- 
    ra_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_403_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(131)); -- 
    -- CP-element group 132:  transition  input  output  no-bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	128 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_403_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Sample/rr
      -- 
    ca_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_403_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(132)); -- 
    rr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(132), ack => ADD_u64_u64_408_inst_req_0); -- 
    -- CP-element group 133:  transition  input  no-bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Sample/ra
      -- 
    ra_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_408_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  no-bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	128 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (27) 
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u64_u64_408_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_offset_calculated
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_resized_0
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_scaled_0
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_computed_0
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_resize_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_resize_0/$exit
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_resize_0/index_resize_req
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_resize_0/index_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_scale_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_scale_0/$exit
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_scale_0/scale_rename_req
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_index_scale_0/scale_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_final_index_sum_regn/$entry
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_final_index_sum_regn/$exit
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_final_index_sum_regn/req
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_final_index_sum_regn/ack
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/array_obj_ref_412_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_request/$entry
      -- CP-element group 134: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_request/req
      -- 
    ca_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_408_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(134)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(134), ack => addr_of_413_final_reg_req_0); -- 
    -- CP-element group 135:  transition  input  no-bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	141 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_request/$exit
      -- CP-element group 135: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_request/ack
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_413_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(135)); -- 
    -- CP-element group 136:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	128 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (24) 
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_complete/$exit
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/addr_of_413_complete/ack
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_address_calculated
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_word_address_calculated
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_root_address_calculated
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_address_resized
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_addr_resize/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_addr_resize/$exit
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_addr_resize/base_resize_req
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_addr_resize/base_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_plus_offset/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_plus_offset/$exit
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_plus_offset/sum_rename_req
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_base_plus_offset/sum_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_word_addrgen/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_word_addrgen/$exit
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_word_addrgen/root_register_req
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_word_addrgen/root_register_ack
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/word_0/rr
      -- 
    ack_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_413_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(136)); -- 
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(136), ack => ptr_deref_417_load_0_req_0); -- 
    -- CP-element group 137:  transition  input  no-bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (5) 
      -- CP-element group 137: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/$exit
      -- CP-element group 137: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/word_0/$exit
      -- CP-element group 137: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Sample/word_access_start/word_0/ra
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_417_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  no-bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	128 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (12) 
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/$exit
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/word_0/$exit
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/word_access_complete/word_0/ca
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/ptr_deref_417_Merge/$entry
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/ptr_deref_417_Merge/$exit
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/ptr_deref_417_Merge/merge_req
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ptr_deref_417_Update/ptr_deref_417_Merge/merge_ack
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Sample/rr
      -- 
    ca_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_417_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(138)); -- 
    rr_1977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(138), ack => ADD_u16_u16_423_inst_req_0); -- 
    -- CP-element group 139:  transition  input  no-bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Sample/ra
      -- 
    ra_1978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_423_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(139)); -- 
    -- CP-element group 140:  transition  input  no-bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	128 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/ADD_u16_u16_423_Update/ca
      -- 
    ca_1983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_423_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(140)); -- 
    -- CP-element group 141:  join  transition  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	135 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	13 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_226/assign_stmt_398_to_assign_stmt_424/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(135) & checkNodeComputeEngine_CP_1062_elements(140);
      gj_checkNodeComputeEngine_cp_element_group_141 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	14 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (7) 
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/$entry
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_update_start_
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Update/cr
      -- 
    rr_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(142), ack => ADD_u16_u16_438_inst_req_0); -- 
    cr_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(142), ack => ADD_u16_u16_438_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(142) <= checkNodeComputeEngine_CP_1062_elements(14);
    -- CP-element group 143:  transition  input  no-bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Sample/ra
      -- 
    ra_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_438_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(143)); -- 
    -- CP-element group 144:  transition  input  no-bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	15 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_226/assign_stmt_439/$exit
      -- CP-element group 144: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_226/assign_stmt_439/ADD_u16_u16_438_Update/ca
      -- 
    ca_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_438_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(144)); -- 
    -- CP-element group 145:  fork  transition  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	16 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	149 
    -- CP-element group 145: 	151 
    -- CP-element group 145: 	153 
    -- CP-element group 145: 	155 
    -- CP-element group 145: 	157 
    -- CP-element group 145:  members (24) 
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_complete/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_complete/req
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/word_0/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/word_0/cr
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_update_start_
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Update/cr
      -- 
    rr_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => ADD_u16_u16_475_inst_req_0); -- 
    cr_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => ADD_u16_u16_475_inst_req_1); -- 
    cr_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => type_cast_479_inst_req_1); -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => addr_of_484_final_reg_req_1); -- 
    cr_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => ptr_deref_488_load_0_req_1); -- 
    cr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => type_cast_492_inst_req_1); -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(145), ack => SLT_f64_u1_498_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(145) <= checkNodeComputeEngine_CP_1062_elements(16);
    -- CP-element group 146:  transition  input  no-bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Sample/ra
      -- 
    ra_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_475_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(146)); -- 
    -- CP-element group 147:  transition  input  output  no-bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ADD_u16_u16_475_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Sample/rr
      -- 
    ca_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_475_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(147)); -- 
    rr_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(147), ack => type_cast_479_inst_req_0); -- 
    -- CP-element group 148:  transition  input  no-bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Sample/ra
      -- 
    ra_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  no-bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	145 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (27) 
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_479_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_root_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_offset_calculated
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_resized_0
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_scaled_0
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_computed_0
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_resize_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_resize_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_resize_0/index_resize_req
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_resize_0/index_resize_ack
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_scale_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_scale_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_scale_0/scale_rename_req
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_index_scale_0/scale_rename_ack
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_final_index_sum_regn/$entry
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_final_index_sum_regn/$exit
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_final_index_sum_regn/req
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_final_index_sum_regn/ack
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_base_plus_offset/$entry
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_base_plus_offset/$exit
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_base_plus_offset/sum_rename_req
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/array_obj_ref_483_base_plus_offset/sum_rename_ack
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_request/$entry
      -- CP-element group 149: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_request/req
      -- 
    ca_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(149)); -- 
    req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(149), ack => addr_of_484_final_reg_req_0); -- 
    -- CP-element group 150:  transition  input  no-bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	158 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_request/$exit
      -- CP-element group 150: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_request/ack
      -- 
    ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_484_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(150)); -- 
    -- CP-element group 151:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	145 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (24) 
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_complete/$exit
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/addr_of_484_complete/ack
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_word_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_root_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_address_resized
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_addr_resize/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_addr_resize/$exit
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_addr_resize/base_resize_req
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_addr_resize/base_resize_ack
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_plus_offset/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_plus_offset/$exit
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_plus_offset/sum_rename_req
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_base_plus_offset/sum_rename_ack
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_word_addrgen/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_word_addrgen/$exit
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_word_addrgen/root_register_req
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_word_addrgen/root_register_ack
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/word_0/$entry
      -- CP-element group 151: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/word_0/rr
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_484_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(151)); -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(151), ack => ptr_deref_488_load_0_req_0); -- 
    -- CP-element group 152:  transition  input  no-bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (5) 
      -- CP-element group 152: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/$exit
      -- CP-element group 152: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/word_0/$exit
      -- CP-element group 152: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Sample/word_access_start/word_0/ra
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_load_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  no-bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	145 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (12) 
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/$exit
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/word_0/$exit
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/word_access_complete/word_0/ca
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/ptr_deref_488_Merge/$entry
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/ptr_deref_488_Merge/$exit
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/ptr_deref_488_Merge/merge_req
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/ptr_deref_488_Update/ptr_deref_488_Merge/merge_ack
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Sample/rr
      -- 
    ca_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_488_load_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(153)); -- 
    rr_2128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(153), ack => type_cast_492_inst_req_0); -- 
    -- CP-element group 154:  transition  input  no-bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Sample/ra
      -- 
    ra_2129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(154)); -- 
    -- CP-element group 155:  transition  input  output  no-bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	145 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/type_cast_492_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Sample/rr
      -- 
    ca_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(155)); -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(155), ack => SLT_f64_u1_498_inst_req_0); -- 
    -- CP-element group 156:  transition  input  no-bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Sample/ra
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_498_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(156)); -- 
    -- CP-element group 157:  transition  input  no-bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	145 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/SLT_f64_u1_498_Update/ca
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_498_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(157)); -- 
    -- CP-element group 158:  join  transition  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	150 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	17 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_226/assign_stmt_476_to_assign_stmt_499/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(150) & checkNodeComputeEngine_CP_1062_elements(157);
      gj_checkNodeComputeEngine_cp_element_group_158 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	17 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_226/if_stmt_500_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(159) <= checkNodeComputeEngine_CP_1062_elements(17);
    -- CP-element group 160:  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	17 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_226/if_stmt_500_eval_test/$entry
      -- CP-element group 160: 	 branch_block_stmt_226/if_stmt_500_eval_test/$exit
      -- CP-element group 160: 	 branch_block_stmt_226/if_stmt_500_eval_test/branch_req
      -- 
    branch_req_2156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(160), ack => if_stmt_500_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(160) <= checkNodeComputeEngine_CP_1062_elements(17);
    -- CP-element group 161:  branch  place  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	164 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_226/R_iNsTr_49_501_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(161) <= checkNodeComputeEngine_CP_1062_elements(160);
    -- CP-element group 162:  transition  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_226/if_stmt_500_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(162) <= checkNodeComputeEngine_CP_1062_elements(161);
    -- CP-element group 163:  transition  input  no-bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_226/if_stmt_500_if_link/$exit
      -- CP-element group 163: 	 branch_block_stmt_226/if_stmt_500_if_link/if_choice_transition
      -- 
    if_choice_transition_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(163)); -- 
    -- CP-element group 164:  transition  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_226/if_stmt_500_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(164) <= checkNodeComputeEngine_CP_1062_elements(161);
    -- CP-element group 165:  transition  input  no-bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_226/if_stmt_500_else_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_226/if_stmt_500_else_link/else_choice_transition
      -- 
    else_choice_transition_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(165)); -- 
    -- CP-element group 166:  place  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	163 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	342 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_226/bb_8_bb_9
      -- 
    checkNodeComputeEngine_CP_1062_elements(166) <= checkNodeComputeEngine_CP_1062_elements(163);
    -- CP-element group 167:  place  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	345 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_226/bb_8_bb_10
      -- 
    checkNodeComputeEngine_CP_1062_elements(167) <= checkNodeComputeEngine_CP_1062_elements(165);
    -- CP-element group 168:  fork  transition  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	18 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (7) 
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/$entry
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_update_start_
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Update/cr
      -- 
    rr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(168), ack => SUB_f32_f32_511_inst_req_0); -- 
    cr_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(168), ack => SUB_f32_f32_511_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(168) <= checkNodeComputeEngine_CP_1062_elements(18);
    -- CP-element group 169:  transition  input  no-bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Sample/ra
      -- 
    ra_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_511_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(169)); -- 
    -- CP-element group 170:  transition  input  no-bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	19 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_226/assign_stmt_512/$exit
      -- CP-element group 170: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_226/assign_stmt_512/SUB_f32_f32_511_Update/ca
      -- 
    ca_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_511_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(170)); -- 
    -- CP-element group 171:  fork  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	20 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (7) 
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/$entry
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_update_start_
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Sample/rr
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Update/cr
      -- 
    rr_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(171), ack => EQ_u16_u1_525_inst_req_0); -- 
    cr_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(171), ack => EQ_u16_u1_525_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(171) <= checkNodeComputeEngine_CP_1062_elements(20);
    -- CP-element group 172:  transition  input  no-bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Sample/ra
      -- 
    ra_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_525_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(172)); -- 
    -- CP-element group 173:  transition  input  no-bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	21 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_226/assign_stmt_526/$exit
      -- CP-element group 173: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_226/assign_stmt_526/EQ_u16_u1_525_Update/ca
      -- 
    ca_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_525_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(173)); -- 
    -- CP-element group 174:  transition  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	21 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_226/if_stmt_527_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(174) <= checkNodeComputeEngine_CP_1062_elements(21);
    -- CP-element group 175:  transition  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	21 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_226/if_stmt_527_eval_test/$entry
      -- CP-element group 175: 	 branch_block_stmt_226/if_stmt_527_eval_test/$exit
      -- CP-element group 175: 	 branch_block_stmt_226/if_stmt_527_eval_test/branch_req
      -- 
    branch_req_2209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(175), ack => if_stmt_527_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(175) <= checkNodeComputeEngine_CP_1062_elements(21);
    -- CP-element group 176:  branch  place  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_226/R_iNsTr_53_528_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(176) <= checkNodeComputeEngine_CP_1062_elements(175);
    -- CP-element group 177:  transition  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_226/if_stmt_527_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(177) <= checkNodeComputeEngine_CP_1062_elements(176);
    -- CP-element group 178:  transition  input  no-bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_226/if_stmt_527_if_link/$exit
      -- CP-element group 178: 	 branch_block_stmt_226/if_stmt_527_if_link/if_choice_transition
      -- 
    if_choice_transition_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_527_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(178)); -- 
    -- CP-element group 179:  transition  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_226/if_stmt_527_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(179) <= checkNodeComputeEngine_CP_1062_elements(176);
    -- CP-element group 180:  transition  input  no-bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_226/if_stmt_527_else_link/$exit
      -- CP-element group 180: 	 branch_block_stmt_226/if_stmt_527_else_link/else_choice_transition
      -- 
    else_choice_transition_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_527_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(180)); -- 
    -- CP-element group 181:  place  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	365 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_226/bb_10_bb_14
      -- 
    checkNodeComputeEngine_CP_1062_elements(181) <= checkNodeComputeEngine_CP_1062_elements(178);
    -- CP-element group 182:  place  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	356 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_226/bb_10_bb_11
      -- 
    checkNodeComputeEngine_CP_1062_elements(182) <= checkNodeComputeEngine_CP_1062_elements(180);
    -- CP-element group 183:  fork  transition  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	22 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	187 
    -- CP-element group 183: 	189 
    -- CP-element group 183: 	190 
    -- CP-element group 183: 	191 
    -- CP-element group 183:  members (19) 
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_update_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_update_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_update_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_update_start_
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Update/cr
      -- 
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => SLT_f64_u1_538_inst_req_0); -- 
    cr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => SLT_f64_u1_538_inst_req_1); -- 
    cr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => type_cast_542_inst_req_1); -- 
    cr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => XOR_u8_u8_547_inst_req_1); -- 
    rr_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => EQ_u8_u1_553_inst_req_0); -- 
    cr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(183), ack => EQ_u8_u1_553_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(183) <= checkNodeComputeEngine_CP_1062_elements(22);
    -- CP-element group 184:  transition  input  no-bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Sample/ra
      -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_538_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  no-bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/SLT_f64_u1_538_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Sample/rr
      -- 
    ca_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_538_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(185)); -- 
    rr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(185), ack => type_cast_542_inst_req_0); -- 
    -- CP-element group 186:  transition  input  no-bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Sample/ra
      -- 
    ra_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  no-bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/type_cast_542_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Sample/rr
      -- 
    ca_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(187)); -- 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(187), ack => XOR_u8_u8_547_inst_req_0); -- 
    -- CP-element group 188:  transition  input  no-bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Sample/ra
      -- 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u8_u8_547_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(188)); -- 
    -- CP-element group 189:  transition  input  no-bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	183 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	192 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/XOR_u8_u8_547_Update/ca
      -- 
    ca_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u8_u8_547_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(189)); -- 
    -- CP-element group 190:  transition  input  no-bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	183 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Sample/ra
      -- 
    ra_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_553_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(190)); -- 
    -- CP-element group 191:  transition  input  no-bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	183 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/EQ_u8_u1_553_Update/ca
      -- 
    ca_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_553_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(191)); -- 
    -- CP-element group 192:  join  transition  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	189 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	23 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_226/assign_stmt_539_to_assign_stmt_554/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(189) & checkNodeComputeEngine_CP_1062_elements(191);
      gj_checkNodeComputeEngine_cp_element_group_192 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  transition  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	23 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_226/if_stmt_555_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(193) <= checkNodeComputeEngine_CP_1062_elements(23);
    -- CP-element group 194:  transition  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	23 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_226/if_stmt_555_eval_test/$entry
      -- CP-element group 194: 	 branch_block_stmt_226/if_stmt_555_eval_test/$exit
      -- CP-element group 194: 	 branch_block_stmt_226/if_stmt_555_eval_test/branch_req
      -- 
    branch_req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(194), ack => if_stmt_555_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(194) <= checkNodeComputeEngine_CP_1062_elements(23);
    -- CP-element group 195:  branch  place  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_226/R_iNsTr_59_556_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(195) <= checkNodeComputeEngine_CP_1062_elements(194);
    -- CP-element group 196:  transition  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_226/if_stmt_555_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(196) <= checkNodeComputeEngine_CP_1062_elements(195);
    -- CP-element group 197:  transition  input  no-bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	200 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_226/if_stmt_555_if_link/$exit
      -- CP-element group 197: 	 branch_block_stmt_226/if_stmt_555_if_link/if_choice_transition
      -- 
    if_choice_transition_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_555_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(197)); -- 
    -- CP-element group 198:  transition  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_226/if_stmt_555_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(198) <= checkNodeComputeEngine_CP_1062_elements(195);
    -- CP-element group 199:  transition  input  no-bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_226/if_stmt_555_else_link/$exit
      -- CP-element group 199: 	 branch_block_stmt_226/if_stmt_555_else_link/else_choice_transition
      -- 
    else_choice_transition_2296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_555_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(199)); -- 
    -- CP-element group 200:  place  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	197 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	376 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_226/bb_11_bb_14
      -- 
    checkNodeComputeEngine_CP_1062_elements(200) <= checkNodeComputeEngine_CP_1062_elements(197);
    -- CP-element group 201:  place  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	359 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_226/bb_11_bb_12
      -- 
    checkNodeComputeEngine_CP_1062_elements(201) <= checkNodeComputeEngine_CP_1062_elements(199);
    -- CP-element group 202:  fork  transition  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	24 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (7) 
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/$entry
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_update_start_
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Sample/rr
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Update/cr
      -- 
    rr_2309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(202), ack => SLT_f32_u1_565_inst_req_0); -- 
    cr_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(202), ack => SLT_f32_u1_565_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(202) <= checkNodeComputeEngine_CP_1062_elements(24);
    -- CP-element group 203:  transition  input  no-bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Sample/ra
      -- 
    ra_2310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_565_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(203)); -- 
    -- CP-element group 204:  transition  input  no-bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	25 
    -- CP-element group 204:  members (4) 
      -- CP-element group 204: 	 branch_block_stmt_226/assign_stmt_566/$exit
      -- CP-element group 204: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_226/assign_stmt_566/SLT_f32_u1_565_Update/ca
      -- 
    ca_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f32_u1_565_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(204)); -- 
    -- CP-element group 205:  transition  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	25 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_226/if_stmt_567_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(205) <= checkNodeComputeEngine_CP_1062_elements(25);
    -- CP-element group 206:  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	25 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_226/if_stmt_567_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_226/if_stmt_567_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_226/if_stmt_567_eval_test/branch_req
      -- 
    branch_req_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(206), ack => if_stmt_567_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(206) <= checkNodeComputeEngine_CP_1062_elements(25);
    -- CP-element group 207:  branch  place  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	210 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_226/R_iNsTr_68_568_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(207) <= checkNodeComputeEngine_CP_1062_elements(206);
    -- CP-element group 208:  transition  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_226/if_stmt_567_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(208) <= checkNodeComputeEngine_CP_1062_elements(207);
    -- CP-element group 209:  transition  input  no-bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	212 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_226/if_stmt_567_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_226/if_stmt_567_if_link/if_choice_transition
      -- 
    if_choice_transition_2328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_567_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(209)); -- 
    -- CP-element group 210:  transition  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	207 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_226/if_stmt_567_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(210) <= checkNodeComputeEngine_CP_1062_elements(207);
    -- CP-element group 211:  transition  input  no-bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_226/if_stmt_567_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_226/if_stmt_567_else_link/else_choice_transition
      -- 
    else_choice_transition_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_567_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(211)); -- 
    -- CP-element group 212:  place  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	209 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	362 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_226/bb_12_bb_13
      -- 
    checkNodeComputeEngine_CP_1062_elements(212) <= checkNodeComputeEngine_CP_1062_elements(209);
    -- CP-element group 213:  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	386 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_226/bb_12_bb_14
      -- 
    checkNodeComputeEngine_CP_1062_elements(213) <= checkNodeComputeEngine_CP_1062_elements(211);
    -- CP-element group 214:  fork  transition  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	27 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214: 	218 
    -- CP-element group 214:  members (10) 
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/$entry
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_update_start_
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_update_start_
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Update/cr
      -- 
    rr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(214), ack => ADD_u16_u16_614_inst_req_0); -- 
    cr_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(214), ack => ADD_u16_u16_614_inst_req_1); -- 
    cr_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(214), ack => EQ_u16_u1_619_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(214) <= checkNodeComputeEngine_CP_1062_elements(27);
    -- CP-element group 215:  transition  input  no-bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Sample/ra
      -- 
    ra_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_614_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(215)); -- 
    -- CP-element group 216:  transition  input  output  no-bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/ADD_u16_u16_614_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Sample/rr
      -- 
    ca_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_614_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(216)); -- 
    rr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(216), ack => EQ_u16_u1_619_inst_req_0); -- 
    -- CP-element group 217:  transition  input  no-bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Sample/ra
      -- 
    ra_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_619_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(217)); -- 
    -- CP-element group 218:  transition  input  no-bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	214 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	28 
    -- CP-element group 218:  members (4) 
      -- CP-element group 218: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/$exit
      -- CP-element group 218: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_226/assign_stmt_615_to_assign_stmt_620/EQ_u16_u1_619_Update/ca
      -- 
    ca_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_619_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(218)); -- 
    -- CP-element group 219:  transition  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	28 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_226/if_stmt_621_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(219) <= checkNodeComputeEngine_CP_1062_elements(28);
    -- CP-element group 220:  transition  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	28 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_226/if_stmt_621_eval_test/$entry
      -- CP-element group 220: 	 branch_block_stmt_226/if_stmt_621_eval_test/$exit
      -- CP-element group 220: 	 branch_block_stmt_226/if_stmt_621_eval_test/branch_req
      -- 
    branch_req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(220), ack => if_stmt_621_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(220) <= checkNodeComputeEngine_CP_1062_elements(28);
    -- CP-element group 221:  branch  place  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221: 	224 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_226/R_exitcond1_622_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(221) <= checkNodeComputeEngine_CP_1062_elements(220);
    -- CP-element group 222:  transition  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 branch_block_stmt_226/if_stmt_621_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(222) <= checkNodeComputeEngine_CP_1062_elements(221);
    -- CP-element group 223:  transition  input  no-bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	226 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_226/if_stmt_621_if_link/$exit
      -- CP-element group 223: 	 branch_block_stmt_226/if_stmt_621_if_link/if_choice_transition
      -- 
    if_choice_transition_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_621_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(223)); -- 
    -- CP-element group 224:  transition  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	221 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_226/if_stmt_621_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(224) <= checkNodeComputeEngine_CP_1062_elements(221);
    -- CP-element group 225:  transition  input  no-bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_226/if_stmt_621_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_226/if_stmt_621_else_link/else_choice_transition
      -- 
    else_choice_transition_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_621_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(225)); -- 
    -- CP-element group 226:  place  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	223 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	412 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge
      -- 
    checkNodeComputeEngine_CP_1062_elements(226) <= checkNodeComputeEngine_CP_1062_elements(223);
    -- CP-element group 227:  place  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	311 
    -- CP-element group 227:  members (1) 
      -- CP-element group 227: 	 branch_block_stmt_226/bb_14_bb_8
      -- 
    checkNodeComputeEngine_CP_1062_elements(227) <= checkNodeComputeEngine_CP_1062_elements(225);
    -- CP-element group 228:  fork  transition  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	29 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228: 	232 
    -- CP-element group 228: 	234 
    -- CP-element group 228: 	235 
    -- CP-element group 228: 	236 
    -- CP-element group 228: 	238 
    -- CP-element group 228: 	241 
    -- CP-element group 228: 	242 
    -- CP-element group 228: 	243 
    -- CP-element group 228: 	245 
    -- CP-element group 228:  members (36) 
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_complete/req
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_complete/req
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_update_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_update_start_
      -- 
    rr_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => EQ_u8_u1_641_inst_req_0); -- 
    cr_2400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => EQ_u8_u1_641_inst_req_1); -- 
    req_2414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => MUX_649_inst_req_1); -- 
    cr_2428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => MUL_f32_f32_654_inst_req_1); -- 
    rr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => type_cast_658_inst_req_0); -- 
    cr_2442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => type_cast_658_inst_req_1); -- 
    req_2481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => addr_of_663_final_reg_req_1); -- 
    cr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => ptr_deref_666_store_0_req_1); -- 
    rr_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => ADD_u16_u16_673_inst_req_0); -- 
    cr_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => ADD_u16_u16_673_inst_req_1); -- 
    cr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(228), ack => EQ_u16_u1_678_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(228) <= checkNodeComputeEngine_CP_1062_elements(29);
    -- CP-element group 229:  transition  input  no-bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Sample/ra
      -- 
    ra_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_641_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(229)); -- 
    -- CP-element group 230:  transition  input  output  no-bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u8_u1_641_Update/ca
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_start/$entry
      -- CP-element group 230: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_start/req
      -- 
    ca_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_641_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(230)); -- 
    req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(230), ack => MUX_649_inst_req_0); -- 
    -- CP-element group 231:  transition  input  no-bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	246 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_start/$exit
      -- CP-element group 231: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_start/ack
      -- 
    ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_649_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  no-bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	228 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_complete/$exit
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUX_649_complete/ack
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Sample/rr
      -- 
    ack_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_649_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(232)); -- 
    rr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(232), ack => MUL_f32_f32_654_inst_req_0); -- 
    -- CP-element group 233:  transition  input  no-bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Sample/ra
      -- 
    ra_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_654_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(233)); -- 
    -- CP-element group 234:  transition  input  no-bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	228 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	239 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/MUL_f32_f32_654_Update/ca
      -- 
    ca_2429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_654_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(234)); -- 
    -- CP-element group 235:  transition  input  no-bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	228 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Sample/ra
      -- CP-element group 235: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_sample_completed_
      -- 
    ra_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(235)); -- 
    -- CP-element group 236:  transition  input  output  no-bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	228 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (27) 
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_scale_0/scale_rename_ack
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_scale_0/$exit
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_base_plus_offset/sum_rename_req
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_scale_0/$entry
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_final_index_sum_regn/$entry
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_resize_0/index_resize_ack
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_resize_0/index_resize_req
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_resized_0
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_offset_calculated
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_root_address_calculated
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_base_plus_offset/$entry
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_scaled_0
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_computed_0
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_resize_0/$entry
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_final_index_sum_regn/req
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_request/req
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_request/$entry
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_scale_0/scale_rename_req
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_final_index_sum_regn/ack
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_Update/ca
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_index_resize_0/$exit
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_final_index_sum_regn/$exit
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_base_plus_offset/$exit
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/array_obj_ref_662_base_plus_offset/sum_rename_ack
      -- CP-element group 236: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/type_cast_658_update_completed_
      -- 
    ca_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(236)); -- 
    req_2476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(236), ack => addr_of_663_final_reg_req_0); -- 
    -- CP-element group 237:  transition  input  no-bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	246 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_request/$exit
      -- CP-element group 237: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_request/ack
      -- 
    ack_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_663_final_reg_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(237)); -- 
    -- CP-element group 238:  fork  transition  input  no-bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	228 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (19) 
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_word_addrgen/root_register_ack
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_word_addrgen/root_register_req
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_word_addrgen/$exit
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_word_addrgen/$entry
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_plus_offset/sum_rename_ack
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_plus_offset/sum_rename_req
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_plus_offset/$exit
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_plus_offset/$entry
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_addr_resize/base_resize_ack
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_addr_resize/base_resize_req
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_addr_resize/$exit
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_addr_resize/$entry
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_address_resized
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_root_address_calculated
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_word_address_calculated
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_base_address_calculated
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_complete/ack
      -- CP-element group 238: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/addr_of_663_complete/$exit
      -- 
    ack_2482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_663_final_reg_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	234 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (9) 
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/word_0/rr
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/word_0/$entry
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/$entry
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/ptr_deref_666_Split/split_ack
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/ptr_deref_666_Split/split_req
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/ptr_deref_666_Split/$exit
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/ptr_deref_666_Split/$entry
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_sample_start_
      -- 
    rr_2520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(239), ack => ptr_deref_666_store_0_req_0); -- 
    checkNodeComputeEngine_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(234) & checkNodeComputeEngine_CP_1062_elements(238);
      gj_checkNodeComputeEngine_cp_element_group_239 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  transition  input  no-bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (5) 
      -- CP-element group 240: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/word_0/ra
      -- CP-element group 240: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/word_0/$exit
      -- CP-element group 240: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/word_access_start/$exit
      -- CP-element group 240: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_sample_completed_
      -- 
    ra_2521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_666_store_0_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(240)); -- 
    -- CP-element group 241:  transition  input  no-bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	228 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	246 
    -- CP-element group 241:  members (5) 
      -- CP-element group 241: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/word_0/ca
      -- CP-element group 241: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/word_0/$exit
      -- CP-element group 241: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/word_access_complete/$exit
      -- CP-element group 241: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ptr_deref_666_update_completed_
      -- 
    ca_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_666_store_0_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(241)); -- 
    -- CP-element group 242:  transition  input  no-bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	228 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_sample_completed_
      -- 
    ra_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_673_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(242)); -- 
    -- CP-element group 243:  transition  input  output  no-bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	228 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/ADD_u16_u16_673_Update/ca
      -- 
    ca_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_673_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(243)); -- 
    rr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(243), ack => EQ_u16_u1_678_inst_req_0); -- 
    -- CP-element group 244:  transition  input  no-bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Sample/ra
      -- CP-element group 244: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_sample_completed_
      -- 
    ra_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_678_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(244)); -- 
    -- CP-element group 245:  transition  input  no-bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	228 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Update/ca
      -- CP-element group 245: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/EQ_u16_u1_678_update_completed_
      -- 
    ca_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_678_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(245)); -- 
    -- CP-element group 246:  join  transition  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	231 
    -- CP-element group 246: 	237 
    -- CP-element group 246: 	241 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	30 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_226/assign_stmt_642_to_assign_stmt_679/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(231) & checkNodeComputeEngine_CP_1062_elements(237) & checkNodeComputeEngine_CP_1062_elements(241) & checkNodeComputeEngine_CP_1062_elements(245);
      gj_checkNodeComputeEngine_cp_element_group_246 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  transition  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	30 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_226/if_stmt_680_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(247) <= checkNodeComputeEngine_CP_1062_elements(30);
    -- CP-element group 248:  transition  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	30 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_226/if_stmt_680_eval_test/branch_req
      -- CP-element group 248: 	 branch_block_stmt_226/if_stmt_680_eval_test/$exit
      -- CP-element group 248: 	 branch_block_stmt_226/if_stmt_680_eval_test/$entry
      -- 
    branch_req_2568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(248), ack => if_stmt_680_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(248) <= checkNodeComputeEngine_CP_1062_elements(30);
    -- CP-element group 249:  branch  place  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (1) 
      -- CP-element group 249: 	 branch_block_stmt_226/R_exitcond_681_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(249) <= checkNodeComputeEngine_CP_1062_elements(248);
    -- CP-element group 250:  transition  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (1) 
      -- CP-element group 250: 	 branch_block_stmt_226/if_stmt_680_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(250) <= checkNodeComputeEngine_CP_1062_elements(249);
    -- CP-element group 251:  transition  input  no-bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	254 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_226/if_stmt_680_if_link/if_choice_transition
      -- CP-element group 251: 	 branch_block_stmt_226/if_stmt_680_if_link/$exit
      -- 
    if_choice_transition_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_680_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(251)); -- 
    -- CP-element group 252:  transition  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (1) 
      -- CP-element group 252: 	 branch_block_stmt_226/if_stmt_680_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(252) <= checkNodeComputeEngine_CP_1062_elements(249);
    -- CP-element group 253:  transition  input  no-bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (2) 
      -- CP-element group 253: 	 branch_block_stmt_226/if_stmt_680_else_link/else_choice_transition
      -- CP-element group 253: 	 branch_block_stmt_226/if_stmt_680_else_link/$exit
      -- 
    else_choice_transition_2577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_680_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(253)); -- 
    -- CP-element group 254:  place  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	251 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	425 
    -- CP-element group 254:  members (1) 
      -- CP-element group 254: 	 branch_block_stmt_226/xx_x_crit_edge_xx_x_crit_edge9x_xloopexit
      -- 
    checkNodeComputeEngine_CP_1062_elements(254) <= checkNodeComputeEngine_CP_1062_elements(251);
    -- CP-element group 255:  place  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	304 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph
      -- 
    checkNodeComputeEngine_CP_1062_elements(255) <= checkNodeComputeEngine_CP_1062_elements(253);
    -- CP-element group 256:  fork  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	32 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (7) 
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Sample/rr
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_update_start_
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/$entry
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Update/cr
      -- 
    rr_2590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(256), ack => ULT_u16_u1_692_inst_req_0); -- 
    cr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(256), ack => ULT_u16_u1_692_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(256) <= checkNodeComputeEngine_CP_1062_elements(32);
    -- CP-element group 257:  transition  input  no-bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Sample/ra
      -- CP-element group 257: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_sample_completed_
      -- 
    ra_2591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u16_u1_692_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(257)); -- 
    -- CP-element group 258:  transition  input  no-bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	33 
    -- CP-element group 258:  members (4) 
      -- CP-element group 258: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_226/assign_stmt_693/$exit
      -- CP-element group 258: 	 branch_block_stmt_226/assign_stmt_693/ULT_u16_u1_692_Update/ca
      -- 
    ca_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u16_u1_692_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(258)); -- 
    -- CP-element group 259:  transition  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	33 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (1) 
      -- CP-element group 259: 	 branch_block_stmt_226/if_stmt_694_dead_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(259) <= checkNodeComputeEngine_CP_1062_elements(33);
    -- CP-element group 260:  transition  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	33 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_226/if_stmt_694_eval_test/$entry
      -- CP-element group 260: 	 branch_block_stmt_226/if_stmt_694_eval_test/$exit
      -- CP-element group 260: 	 branch_block_stmt_226/if_stmt_694_eval_test/branch_req
      -- 
    branch_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(260), ack => if_stmt_694_branch_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(260) <= checkNodeComputeEngine_CP_1062_elements(33);
    -- CP-element group 261:  branch  place  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: 	264 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_226/R_iNsTr_33_695_place
      -- 
    checkNodeComputeEngine_CP_1062_elements(261) <= checkNodeComputeEngine_CP_1062_elements(260);
    -- CP-element group 262:  transition  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_226/if_stmt_694_if_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(262) <= checkNodeComputeEngine_CP_1062_elements(261);
    -- CP-element group 263:  transition  input  no-bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	266 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_226/if_stmt_694_if_link/$exit
      -- CP-element group 263: 	 branch_block_stmt_226/if_stmt_694_if_link/if_choice_transition
      -- 
    if_choice_transition_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_694_branch_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(263)); -- 
    -- CP-element group 264:  transition  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	261 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (1) 
      -- CP-element group 264: 	 branch_block_stmt_226/if_stmt_694_else_link/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(264) <= checkNodeComputeEngine_CP_1062_elements(261);
    -- CP-element group 265:  transition  input  no-bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (2) 
      -- CP-element group 265: 	 branch_block_stmt_226/if_stmt_694_else_link/$exit
      -- CP-element group 265: 	 branch_block_stmt_226/if_stmt_694_else_link/else_choice_transition
      -- 
    else_choice_transition_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_694_branch_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(265)); -- 
    -- CP-element group 266:  place  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	263 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	274 
    -- CP-element group 266:  members (1) 
      -- CP-element group 266: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11
      -- 
    checkNodeComputeEngine_CP_1062_elements(266) <= checkNodeComputeEngine_CP_1062_elements(263);
    -- CP-element group 267:  place  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	432 
    -- CP-element group 267:  members (1) 
      -- CP-element group 267: 	 branch_block_stmt_226/xx_x_crit_edge9_xx_x_crit_edge12x_xloopexit
      -- 
    checkNodeComputeEngine_CP_1062_elements(267) <= checkNodeComputeEngine_CP_1062_elements(265);
    -- CP-element group 268:  transition  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	50 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (2) 
      -- CP-element group 268: 	 branch_block_stmt_226/bb_0_bbx_xnph11x_xpreheader_PhiReq/$entry
      -- CP-element group 268: 	 branch_block_stmt_226/bb_0_bbx_xnph11x_xpreheader_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(268) <= checkNodeComputeEngine_CP_1062_elements(50);
    -- CP-element group 269:  place  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (1) 
      -- CP-element group 269: 	 branch_block_stmt_226/merge_stmt_242_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(269) <= checkNodeComputeEngine_CP_1062_elements(268);
    -- CP-element group 270:  transition  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	3 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_226/merge_stmt_242_PhiAck/$entry
      -- CP-element group 270: 	 branch_block_stmt_226/merge_stmt_242_PhiAck/$exit
      -- CP-element group 270: 	 branch_block_stmt_226/merge_stmt_242_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(270) <= checkNodeComputeEngine_CP_1062_elements(269);
    -- CP-element group 271:  transition  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	3 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/$entry
      -- CP-element group 271: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/$entry
      -- CP-element group 271: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(271) <= checkNodeComputeEngine_CP_1062_elements(3);
    -- CP-element group 272:  transition  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (1) 
      -- CP-element group 272: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_251_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(272) is a control-delay.
    cp_element_272_delay: control_delay_element  generic map(name => " 272_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(271), ack => checkNodeComputeEngine_CP_1062_elements(272), clk => clk, reset =>reset);
    -- CP-element group 273:  transition  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	278 
    -- CP-element group 273:  members (4) 
      -- CP-element group 273: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/$exit
      -- CP-element group 273: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/$exit
      -- CP-element group 273: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/$exit
      -- CP-element group 273: 	 branch_block_stmt_226/bbx_xnph11x_xpreheader_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_req
      -- 
    phi_stmt_245_req_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_245_req_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(273), ack => phi_stmt_245_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(273) <= checkNodeComputeEngine_CP_1062_elements(272);
    -- CP-element group 274:  fork  transition  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	266 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (9) 
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Update/cr
      -- 
    rr_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(274), ack => type_cast_248_inst_req_0); -- 
    cr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(274), ack => type_cast_248_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(274) <= checkNodeComputeEngine_CP_1062_elements(266);
    -- CP-element group 275:  transition  input  no-bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (2) 
      -- CP-element group 275: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Sample/ra
      -- 
    ra_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_248_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(275)); -- 
    -- CP-element group 276:  transition  input  no-bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/Update/ca
      -- 
    ca_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_248_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/$exit
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/$exit
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/$exit
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/$exit
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_sources/type_cast_248/SplitProtocol/$exit
      -- CP-element group 277: 	 branch_block_stmt_226/xx_x_crit_edge9_bbx_xnph11_PhiReq/phi_stmt_245/phi_stmt_245_req
      -- 
    phi_stmt_245_req_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_245_req_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(277), ack => phi_stmt_245_req_0); -- 
    checkNodeComputeEngine_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(275) & checkNodeComputeEngine_CP_1062_elements(276);
      gj_checkNodeComputeEngine_cp_element_group_277 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  merge  place  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	273 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (1) 
      -- CP-element group 278: 	 branch_block_stmt_226/merge_stmt_244_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(278) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(273) & checkNodeComputeEngine_CP_1062_elements(277));
    -- CP-element group 279:  transition  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (1) 
      -- CP-element group 279: 	 branch_block_stmt_226/merge_stmt_244_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(279) <= checkNodeComputeEngine_CP_1062_elements(278);
    -- CP-element group 280:  transition  input  no-bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	4 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_226/merge_stmt_244_PhiAck/$exit
      -- CP-element group 280: 	 branch_block_stmt_226/merge_stmt_244_PhiAck/phi_stmt_245_ack
      -- 
    phi_stmt_245_ack_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_245_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(280)); -- 
    -- CP-element group 281:  transition  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	87 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_226/bbx_xnph11_bb_4_PhiReq/$entry
      -- CP-element group 281: 	 branch_block_stmt_226/bbx_xnph11_bb_4_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(281) <= checkNodeComputeEngine_CP_1062_elements(87);
    -- CP-element group 282:  place  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_226/merge_stmt_316_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(282) <= checkNodeComputeEngine_CP_1062_elements(281);
    -- CP-element group 283:  transition  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	6 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_226/merge_stmt_316_PhiAck/$entry
      -- CP-element group 283: 	 branch_block_stmt_226/merge_stmt_316_PhiAck/$exit
      -- CP-element group 283: 	 branch_block_stmt_226/merge_stmt_316_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(283) <= checkNodeComputeEngine_CP_1062_elements(282);
    -- CP-element group 284:  transition  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	86 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_226/bbx_xnph11_bb_3_PhiReq/$entry
      -- CP-element group 284: 	 branch_block_stmt_226/bbx_xnph11_bb_3_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(284) <= checkNodeComputeEngine_CP_1062_elements(86);
    -- CP-element group 285:  place  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_226/merge_stmt_352_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(285) <= checkNodeComputeEngine_CP_1062_elements(284);
    -- CP-element group 286:  transition  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	8 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_226/merge_stmt_352_PhiAck/$entry
      -- CP-element group 286: 	 branch_block_stmt_226/merge_stmt_352_PhiAck/$exit
      -- CP-element group 286: 	 branch_block_stmt_226/merge_stmt_352_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(286) <= checkNodeComputeEngine_CP_1062_elements(285);
    -- CP-element group 287:  fork  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	9 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (9) 
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Update/cr
      -- 
    rr_2708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(287), ack => type_cast_378_inst_req_0); -- 
    cr_2713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(287), ack => type_cast_378_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(287) <= checkNodeComputeEngine_CP_1062_elements(9);
    -- CP-element group 288:  transition  input  no-bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Sample/ra
      -- 
    ra_2709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(288)); -- 
    -- CP-element group 289:  transition  input  no-bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/Update/ca
      -- 
    ca_2714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	295 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/$exit
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/$exit
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/$exit
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_378/SplitProtocol/$exit
      -- CP-element group 290: 	 branch_block_stmt_226/bb_3_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_req
      -- 
    phi_stmt_375_req_2715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_375_req_2715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(290), ack => phi_stmt_375_req_0); -- 
    checkNodeComputeEngine_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(288) & checkNodeComputeEngine_CP_1062_elements(289);
      gj_checkNodeComputeEngine_cp_element_group_290 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	7 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (9) 
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Sample/rr
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Update/cr
      -- 
    rr_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(291), ack => type_cast_380_inst_req_0); -- 
    cr_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(291), ack => type_cast_380_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(291) <= checkNodeComputeEngine_CP_1062_elements(7);
    -- CP-element group 292:  transition  input  no-bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Sample/ra
      -- 
    ra_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(292)); -- 
    -- CP-element group 293:  transition  input  no-bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (2) 
      -- CP-element group 293: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/Update/ca
      -- 
    ca_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/$exit
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/$exit
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/$exit
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/$exit
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_sources/type_cast_380/SplitProtocol/$exit
      -- CP-element group 294: 	 branch_block_stmt_226/bb_4_bb_5_PhiReq/phi_stmt_375/phi_stmt_375_req
      -- 
    phi_stmt_375_req_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_375_req_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(294), ack => phi_stmt_375_req_1); -- 
    checkNodeComputeEngine_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(292) & checkNodeComputeEngine_CP_1062_elements(293);
      gj_checkNodeComputeEngine_cp_element_group_294 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  merge  place  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	290 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (1) 
      -- CP-element group 295: 	 branch_block_stmt_226/merge_stmt_374_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(295) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(290) & checkNodeComputeEngine_CP_1062_elements(294));
    -- CP-element group 296:  transition  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_226/merge_stmt_374_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(296) <= checkNodeComputeEngine_CP_1062_elements(295);
    -- CP-element group 297:  transition  input  no-bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	10 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_226/merge_stmt_374_PhiAck/$exit
      -- CP-element group 297: 	 branch_block_stmt_226/merge_stmt_374_PhiAck/phi_stmt_375_ack
      -- 
    phi_stmt_375_ack_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_375_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(297)); -- 
    -- CP-element group 298:  transition  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	127 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_226/bb_5_bbx_xnph8_PhiReq/$entry
      -- CP-element group 298: 	 branch_block_stmt_226/bb_5_bbx_xnph8_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(298) <= checkNodeComputeEngine_CP_1062_elements(127);
    -- CP-element group 299:  place  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (1) 
      -- CP-element group 299: 	 branch_block_stmt_226/merge_stmt_394_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(299) <= checkNodeComputeEngine_CP_1062_elements(298);
    -- CP-element group 300:  transition  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	12 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_226/merge_stmt_394_PhiAck/$entry
      -- CP-element group 300: 	 branch_block_stmt_226/merge_stmt_394_PhiAck/$exit
      -- CP-element group 300: 	 branch_block_stmt_226/merge_stmt_394_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(300) <= checkNodeComputeEngine_CP_1062_elements(299);
    -- CP-element group 301:  transition  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	13 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/$entry
      -- CP-element group 301: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/$entry
      -- CP-element group 301: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(301) <= checkNodeComputeEngine_CP_1062_elements(13);
    -- CP-element group 302:  transition  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (1) 
      -- CP-element group 302: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_431_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(302) is a control-delay.
    cp_element_302_delay: control_delay_element  generic map(name => " 302_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(301), ack => checkNodeComputeEngine_CP_1062_elements(302), clk => clk, reset =>reset);
    -- CP-element group 303:  transition  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	308 
    -- CP-element group 303:  members (4) 
      -- CP-element group 303: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/$exit
      -- CP-element group 303: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/$exit
      -- CP-element group 303: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/$exit
      -- CP-element group 303: 	 branch_block_stmt_226/bbx_xnph8_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_req
      -- 
    phi_stmt_427_req_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_427_req_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(303), ack => phi_stmt_427_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(303) <= checkNodeComputeEngine_CP_1062_elements(302);
    -- CP-element group 304:  fork  transition  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	255 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (9) 
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Sample/rr
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Update/cr
      -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(304), ack => type_cast_433_inst_req_0); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(304), ack => type_cast_433_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(304) <= checkNodeComputeEngine_CP_1062_elements(255);
    -- CP-element group 305:  transition  input  no-bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Sample/ra
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_433_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(305)); -- 
    -- CP-element group 306:  transition  input  no-bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_433_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/$exit
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/$exit
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/$exit
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_sources/type_cast_433/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_226/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_427/phi_stmt_427_req
      -- 
    phi_stmt_427_req_2795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_427_req_2795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(307), ack => phi_stmt_427_req_1); -- 
    checkNodeComputeEngine_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(305) & checkNodeComputeEngine_CP_1062_elements(306);
      gj_checkNodeComputeEngine_cp_element_group_307 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  merge  place  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	303 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (1) 
      -- CP-element group 308: 	 branch_block_stmt_226/merge_stmt_426_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(308) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(303) & checkNodeComputeEngine_CP_1062_elements(307));
    -- CP-element group 309:  transition  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (1) 
      -- CP-element group 309: 	 branch_block_stmt_226/merge_stmt_426_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(309) <= checkNodeComputeEngine_CP_1062_elements(308);
    -- CP-element group 310:  transition  input  no-bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	14 
    -- CP-element group 310:  members (2) 
      -- CP-element group 310: 	 branch_block_stmt_226/merge_stmt_426_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_226/merge_stmt_426_PhiAck/phi_stmt_427_ack
      -- 
    phi_stmt_427_ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_427_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(310)); -- 
    -- CP-element group 311:  fork  transition  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	227 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311: 	313 
    -- CP-element group 311: 	315 
    -- CP-element group 311: 	316 
    -- CP-element group 311: 	318 
    -- CP-element group 311: 	319 
    -- CP-element group 311: 	321 
    -- CP-element group 311: 	322 
    -- CP-element group 311:  members (33) 
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Sample/rr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Update/cr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/rr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/cr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Sample/rr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Update/cr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Sample/rr
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Update/cr
      -- 
    rr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_449_inst_req_0); -- 
    cr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_449_inst_req_1); -- 
    rr_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_456_inst_req_0); -- 
    cr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_456_inst_req_1); -- 
    rr_2865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_463_inst_req_0); -- 
    cr_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_463_inst_req_1); -- 
    rr_2888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_470_inst_req_0); -- 
    cr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(311), ack => type_cast_470_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(311) <= checkNodeComputeEngine_CP_1062_elements(227);
    -- CP-element group 312:  transition  input  no-bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Sample/ra
      -- 
    ra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_449_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(312)); -- 
    -- CP-element group 313:  transition  input  no-bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (2) 
      -- CP-element group 313: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/Update/ca
      -- 
    ca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_449_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	324 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/$exit
      -- CP-element group 314: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/$exit
      -- CP-element group 314: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_449/SplitProtocol/$exit
      -- CP-element group 314: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_req
      -- 
    phi_stmt_442_req_2826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_442_req_2826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(314), ack => phi_stmt_442_req_1); -- 
    checkNodeComputeEngine_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(312) & checkNodeComputeEngine_CP_1062_elements(313);
      gj_checkNodeComputeEngine_cp_element_group_314 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  transition  input  no-bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	311 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/ra
      -- 
    ra_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(315)); -- 
    -- CP-element group 316:  transition  input  no-bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	311 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/ca
      -- 
    ca_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	324 
    -- CP-element group 317:  members (5) 
      -- CP-element group 317: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/$exit
      -- CP-element group 317: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/$exit
      -- CP-element group 317: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/$exit
      -- CP-element group 317: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/$exit
      -- CP-element group 317: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_req
      -- 
    phi_stmt_450_req_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_450_req_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(317), ack => phi_stmt_450_req_1); -- 
    checkNodeComputeEngine_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(315) & checkNodeComputeEngine_CP_1062_elements(316);
      gj_checkNodeComputeEngine_cp_element_group_317 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  no-bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	311 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Sample/ra
      -- 
    ra_2866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_463_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(318)); -- 
    -- CP-element group 319:  transition  input  no-bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	311 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/Update/ca
      -- 
    ca_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_463_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(319)); -- 
    -- CP-element group 320:  join  transition  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	324 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/$exit
      -- CP-element group 320: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/$exit
      -- CP-element group 320: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/$exit
      -- CP-element group 320: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_463/SplitProtocol/$exit
      -- CP-element group 320: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_req
      -- 
    phi_stmt_457_req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_457_req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(320), ack => phi_stmt_457_req_1); -- 
    checkNodeComputeEngine_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(318) & checkNodeComputeEngine_CP_1062_elements(319);
      gj_checkNodeComputeEngine_cp_element_group_320 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  transition  input  no-bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	311 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Sample/ra
      -- 
    ra_2889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(321)); -- 
    -- CP-element group 322:  transition  input  no-bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	311 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/Update/ca
      -- 
    ca_2894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/$exit
      -- CP-element group 323: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/$exit
      -- CP-element group 323: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/$exit
      -- CP-element group 323: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_470/SplitProtocol/$exit
      -- CP-element group 323: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_req
      -- 
    phi_stmt_464_req_2895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_464_req_2895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(323), ack => phi_stmt_464_req_1); -- 
    checkNodeComputeEngine_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(321) & checkNodeComputeEngine_CP_1062_elements(322);
      gj_checkNodeComputeEngine_cp_element_group_323 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  join  transition  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	314 
    -- CP-element group 324: 	317 
    -- CP-element group 324: 	320 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	335 
    -- CP-element group 324:  members (1) 
      -- CP-element group 324: 	 branch_block_stmt_226/bb_14_bb_8_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(314) & checkNodeComputeEngine_CP_1062_elements(317) & checkNodeComputeEngine_CP_1062_elements(320) & checkNodeComputeEngine_CP_1062_elements(323);
      gj_checkNodeComputeEngine_cp_element_group_324 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  fork  transition  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	15 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325: 	328 
    -- CP-element group 325: 	330 
    -- CP-element group 325: 	332 
    -- CP-element group 325:  members (9) 
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/$entry
      -- CP-element group 325: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(325) <= checkNodeComputeEngine_CP_1062_elements(15);
    -- CP-element group 326:  transition  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/type_cast_447_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(326) is a control-delay.
    cp_element_326_delay: control_delay_element  generic map(name => " 326_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(325), ack => checkNodeComputeEngine_CP_1062_elements(326), clk => clk, reset =>reset);
    -- CP-element group 327:  transition  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	334 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/$exit
      -- CP-element group 327: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_442/phi_stmt_442_req
      -- 
    phi_stmt_442_req_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_442_req_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(327), ack => phi_stmt_442_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(327) <= checkNodeComputeEngine_CP_1062_elements(326);
    -- CP-element group 328:  transition  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	325 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_454_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(328) is a control-delay.
    cp_element_328_delay: control_delay_element  generic map(name => " 328_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(325), ack => checkNodeComputeEngine_CP_1062_elements(328), clk => clk, reset =>reset);
    -- CP-element group 329:  transition  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	334 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/$exit
      -- CP-element group 329: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_sources/$exit
      -- CP-element group 329: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_450/phi_stmt_450_req
      -- 
    phi_stmt_450_req_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_450_req_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(329), ack => phi_stmt_450_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(329) <= checkNodeComputeEngine_CP_1062_elements(328);
    -- CP-element group 330:  transition  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	325 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/type_cast_461_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(330) is a control-delay.
    cp_element_330_delay: control_delay_element  generic map(name => " 330_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(325), ack => checkNodeComputeEngine_CP_1062_elements(330), clk => clk, reset =>reset);
    -- CP-element group 331:  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	334 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/$exit
      -- CP-element group 331: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_sources/$exit
      -- CP-element group 331: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_457/phi_stmt_457_req
      -- 
    phi_stmt_457_req_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_457_req_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(331), ack => phi_stmt_457_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(331) <= checkNodeComputeEngine_CP_1062_elements(330);
    -- CP-element group 332:  transition  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	325 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (1) 
      -- CP-element group 332: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/type_cast_468_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(332) is a control-delay.
    cp_element_332_delay: control_delay_element  generic map(name => " 332_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(325), ack => checkNodeComputeEngine_CP_1062_elements(332), clk => clk, reset =>reset);
    -- CP-element group 333:  transition  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/$exit
      -- CP-element group 333: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_sources/$exit
      -- CP-element group 333: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/phi_stmt_464/phi_stmt_464_req
      -- 
    phi_stmt_464_req_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_464_req_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(333), ack => phi_stmt_464_req_0); -- 
    checkNodeComputeEngine_CP_1062_elements(333) <= checkNodeComputeEngine_CP_1062_elements(332);
    -- CP-element group 334:  join  transition  no-bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	327 
    -- CP-element group 334: 	329 
    -- CP-element group 334: 	331 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (1) 
      -- CP-element group 334: 	 branch_block_stmt_226/bbx_xnph_bb_8_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(327) & checkNodeComputeEngine_CP_1062_elements(329) & checkNodeComputeEngine_CP_1062_elements(331) & checkNodeComputeEngine_CP_1062_elements(333);
      gj_checkNodeComputeEngine_cp_element_group_334 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  merge  place  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	324 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (1) 
      -- CP-element group 335: 	 branch_block_stmt_226/merge_stmt_441_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(335) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(324) & checkNodeComputeEngine_CP_1062_elements(334));
    -- CP-element group 336:  fork  transition  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	338 
    -- CP-element group 336: 	339 
    -- CP-element group 336: 	340 
    -- CP-element group 336:  members (1) 
      -- CP-element group 336: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(336) <= checkNodeComputeEngine_CP_1062_elements(335);
    -- CP-element group 337:  transition  input  no-bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	341 
    -- CP-element group 337:  members (1) 
      -- CP-element group 337: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/phi_stmt_442_ack
      -- 
    phi_stmt_442_ack_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_442_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(337)); -- 
    -- CP-element group 338:  transition  input  no-bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	341 
    -- CP-element group 338:  members (1) 
      -- CP-element group 338: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/phi_stmt_450_ack
      -- 
    phi_stmt_450_ack_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_450_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(338)); -- 
    -- CP-element group 339:  transition  input  no-bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	336 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (1) 
      -- CP-element group 339: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/phi_stmt_457_ack
      -- 
    phi_stmt_457_ack_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_457_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(339)); -- 
    -- CP-element group 340:  transition  input  no-bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	336 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (1) 
      -- CP-element group 340: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/phi_stmt_464_ack
      -- 
    phi_stmt_464_ack_2938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_464_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(340)); -- 
    -- CP-element group 341:  join  transition  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	337 
    -- CP-element group 341: 	338 
    -- CP-element group 341: 	339 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	16 
    -- CP-element group 341:  members (1) 
      -- CP-element group 341: 	 branch_block_stmt_226/merge_stmt_441_PhiAck/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(337) & checkNodeComputeEngine_CP_1062_elements(338) & checkNodeComputeEngine_CP_1062_elements(339) & checkNodeComputeEngine_CP_1062_elements(340);
      gj_checkNodeComputeEngine_cp_element_group_341 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  transition  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	166 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (2) 
      -- CP-element group 342: 	 branch_block_stmt_226/bb_8_bb_9_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_226/bb_8_bb_9_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(342) <= checkNodeComputeEngine_CP_1062_elements(166);
    -- CP-element group 343:  place  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (1) 
      -- CP-element group 343: 	 branch_block_stmt_226/merge_stmt_506_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(343) <= checkNodeComputeEngine_CP_1062_elements(342);
    -- CP-element group 344:  transition  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	18 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_226/merge_stmt_506_PhiAck/$entry
      -- CP-element group 344: 	 branch_block_stmt_226/merge_stmt_506_PhiAck/$exit
      -- CP-element group 344: 	 branch_block_stmt_226/merge_stmt_506_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(344) <= checkNodeComputeEngine_CP_1062_elements(343);
    -- CP-element group 345:  fork  transition  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	167 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (9) 
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Sample/rr
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Update/cr
      -- 
    rr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(345), ack => type_cast_520_inst_req_0); -- 
    cr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(345), ack => type_cast_520_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(345) <= checkNodeComputeEngine_CP_1062_elements(167);
    -- CP-element group 346:  transition  input  no-bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Sample/ra
      -- 
    ra_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(346)); -- 
    -- CP-element group 347:  transition  input  no-bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/Update/ca
      -- 
    ca_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	353 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/$exit
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/$exit
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/$exit
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_520/SplitProtocol/$exit
      -- CP-element group 348: 	 branch_block_stmt_226/bb_8_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_req
      -- 
    phi_stmt_515_req_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_515_req_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(348), ack => phi_stmt_515_req_1); -- 
    checkNodeComputeEngine_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(346) & checkNodeComputeEngine_CP_1062_elements(347);
      gj_checkNodeComputeEngine_cp_element_group_348 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	19 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (9) 
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Sample/rr
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Update/cr
      -- 
    rr_2995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(349), ack => type_cast_518_inst_req_0); -- 
    cr_3000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(349), ack => type_cast_518_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(349) <= checkNodeComputeEngine_CP_1062_elements(19);
    -- CP-element group 350:  transition  input  no-bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Sample/ra
      -- 
    ra_2996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(350)); -- 
    -- CP-element group 351:  transition  input  no-bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (2) 
      -- CP-element group 351: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/Update/ca
      -- 
    ca_3001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(351)); -- 
    -- CP-element group 352:  join  transition  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/$exit
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/$exit
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/$exit
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/$exit
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_sources/type_cast_518/SplitProtocol/$exit
      -- CP-element group 352: 	 branch_block_stmt_226/bb_9_bb_10_PhiReq/phi_stmt_515/phi_stmt_515_req
      -- 
    phi_stmt_515_req_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_515_req_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(352), ack => phi_stmt_515_req_0); -- 
    checkNodeComputeEngine_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(350) & checkNodeComputeEngine_CP_1062_elements(351);
      gj_checkNodeComputeEngine_cp_element_group_352 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  merge  place  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	348 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (1) 
      -- CP-element group 353: 	 branch_block_stmt_226/merge_stmt_514_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(353) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(348) & checkNodeComputeEngine_CP_1062_elements(352));
    -- CP-element group 354:  transition  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (1) 
      -- CP-element group 354: 	 branch_block_stmt_226/merge_stmt_514_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(354) <= checkNodeComputeEngine_CP_1062_elements(353);
    -- CP-element group 355:  transition  input  no-bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	20 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_226/merge_stmt_514_PhiAck/$exit
      -- CP-element group 355: 	 branch_block_stmt_226/merge_stmt_514_PhiAck/phi_stmt_515_ack
      -- 
    phi_stmt_515_ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_515_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(355)); -- 
    -- CP-element group 356:  transition  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	182 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (2) 
      -- CP-element group 356: 	 branch_block_stmt_226/bb_10_bb_11_PhiReq/$entry
      -- CP-element group 356: 	 branch_block_stmt_226/bb_10_bb_11_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(356) <= checkNodeComputeEngine_CP_1062_elements(182);
    -- CP-element group 357:  place  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (1) 
      -- CP-element group 357: 	 branch_block_stmt_226/merge_stmt_533_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(357) <= checkNodeComputeEngine_CP_1062_elements(356);
    -- CP-element group 358:  transition  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	22 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_226/merge_stmt_533_PhiAck/$entry
      -- CP-element group 358: 	 branch_block_stmt_226/merge_stmt_533_PhiAck/$exit
      -- CP-element group 358: 	 branch_block_stmt_226/merge_stmt_533_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(358) <= checkNodeComputeEngine_CP_1062_elements(357);
    -- CP-element group 359:  transition  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	201 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (2) 
      -- CP-element group 359: 	 branch_block_stmt_226/bb_11_bb_12_PhiReq/$entry
      -- CP-element group 359: 	 branch_block_stmt_226/bb_11_bb_12_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(359) <= checkNodeComputeEngine_CP_1062_elements(201);
    -- CP-element group 360:  place  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (1) 
      -- CP-element group 360: 	 branch_block_stmt_226/merge_stmt_561_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(360) <= checkNodeComputeEngine_CP_1062_elements(359);
    -- CP-element group 361:  transition  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	24 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_226/merge_stmt_561_PhiAck/$entry
      -- CP-element group 361: 	 branch_block_stmt_226/merge_stmt_561_PhiAck/$exit
      -- CP-element group 361: 	 branch_block_stmt_226/merge_stmt_561_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(361) <= checkNodeComputeEngine_CP_1062_elements(360);
    -- CP-element group 362:  transition  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	212 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_226/bb_12_bb_13_PhiReq/$entry
      -- CP-element group 362: 	 branch_block_stmt_226/bb_12_bb_13_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(362) <= checkNodeComputeEngine_CP_1062_elements(212);
    -- CP-element group 363:  place  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (1) 
      -- CP-element group 363: 	 branch_block_stmt_226/merge_stmt_573_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(363) <= checkNodeComputeEngine_CP_1062_elements(362);
    -- CP-element group 364:  transition  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	26 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_226/merge_stmt_573_PhiAck/$entry
      -- CP-element group 364: 	 branch_block_stmt_226/merge_stmt_573_PhiAck/$exit
      -- CP-element group 364: 	 branch_block_stmt_226/merge_stmt_573_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(364) <= checkNodeComputeEngine_CP_1062_elements(363);
    -- CP-element group 365:  fork  transition  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	181 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: 	367 
    -- CP-element group 365: 	369 
    -- CP-element group 365: 	370 
    -- CP-element group 365: 	372 
    -- CP-element group 365: 	373 
    -- CP-element group 365:  members (25) 
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Update/cr
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Update/cr
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Update/cr
      -- 
    rr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_579_inst_req_0); -- 
    cr_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_579_inst_req_1); -- 
    rr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_592_inst_req_0); -- 
    cr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_592_inst_req_1); -- 
    rr_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_602_inst_req_0); -- 
    cr_3113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(365), ack => type_cast_602_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(365) <= checkNodeComputeEngine_CP_1062_elements(181);
    -- CP-element group 366:  transition  input  no-bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (2) 
      -- CP-element group 366: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Sample/ra
      -- 
    ra_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(366)); -- 
    -- CP-element group 367:  transition  input  no-bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/Update/ca
      -- 
    ca_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(367)); -- 
    -- CP-element group 368:  join  transition  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	375 
    -- CP-element group 368:  members (5) 
      -- CP-element group 368: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/$exit
      -- CP-element group 368: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$exit
      -- CP-element group 368: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/$exit
      -- CP-element group 368: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_579/SplitProtocol/$exit
      -- CP-element group 368: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_req
      -- 
    phi_stmt_576_req_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_576_req_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(368), ack => phi_stmt_576_req_0); -- 
    checkNodeComputeEngine_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(366) & checkNodeComputeEngine_CP_1062_elements(367);
      gj_checkNodeComputeEngine_cp_element_group_368 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  transition  input  no-bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Sample/ra
      -- 
    ra_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(369)); -- 
    -- CP-element group 370:  transition  input  no-bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/Update/ca
      -- 
    ca_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	375 
    -- CP-element group 371:  members (5) 
      -- CP-element group 371: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/$exit
      -- CP-element group 371: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- CP-element group 371: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/$exit
      -- CP-element group 371: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_592/SplitProtocol/$exit
      -- CP-element group 371: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    phi_stmt_589_req_3092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_req_3092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(371), ack => phi_stmt_589_req_0); -- 
    checkNodeComputeEngine_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(369) & checkNodeComputeEngine_CP_1062_elements(370);
      gj_checkNodeComputeEngine_cp_element_group_371 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  transition  input  no-bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	365 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (2) 
      -- CP-element group 372: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Sample/ra
      -- 
    ra_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(372)); -- 
    -- CP-element group 373:  transition  input  no-bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	365 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (2) 
      -- CP-element group 373: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/Update/ca
      -- 
    ca_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_602_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/$exit
      -- CP-element group 374: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$exit
      -- CP-element group 374: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/$exit
      -- CP-element group 374: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_602/SplitProtocol/$exit
      -- CP-element group 374: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_req
      -- 
    phi_stmt_599_req_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_599_req_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(374), ack => phi_stmt_599_req_0); -- 
    checkNodeComputeEngine_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(372) & checkNodeComputeEngine_CP_1062_elements(373);
      gj_checkNodeComputeEngine_cp_element_group_374 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  join  transition  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	368 
    -- CP-element group 375: 	371 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	406 
    -- CP-element group 375:  members (1) 
      -- CP-element group 375: 	 branch_block_stmt_226/bb_10_bb_14_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(368) & checkNodeComputeEngine_CP_1062_elements(371) & checkNodeComputeEngine_CP_1062_elements(374);
      gj_checkNodeComputeEngine_cp_element_group_375 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  fork  transition  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	200 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376: 	379 
    -- CP-element group 376: 	380 
    -- CP-element group 376: 	382 
    -- CP-element group 376: 	383 
    -- CP-element group 376:  members (19) 
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Sample/rr
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Update/cr
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Sample/rr
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Update/cr
      -- 
    rr_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(376), ack => type_cast_594_inst_req_0); -- 
    cr_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(376), ack => type_cast_594_inst_req_1); -- 
    rr_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(376), ack => type_cast_604_inst_req_0); -- 
    cr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(376), ack => type_cast_604_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(376) <= checkNodeComputeEngine_CP_1062_elements(200);
    -- CP-element group 377:  transition  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_582_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(377) is a control-delay.
    cp_element_377_delay: control_delay_element  generic map(name => " 377_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(376), ack => checkNodeComputeEngine_CP_1062_elements(377), clk => clk, reset =>reset);
    -- CP-element group 378:  transition  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	385 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/$exit
      -- CP-element group 378: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$exit
      -- CP-element group 378: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_req
      -- 
    phi_stmt_576_req_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_576_req_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(378), ack => phi_stmt_576_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(378) <= checkNodeComputeEngine_CP_1062_elements(377);
    -- CP-element group 379:  transition  input  no-bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	376 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (2) 
      -- CP-element group 379: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Sample/ra
      -- 
    ra_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(379)); -- 
    -- CP-element group 380:  transition  input  no-bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	376 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/Update/ca
      -- 
    ca_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(380)); -- 
    -- CP-element group 381:  join  transition  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	385 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/$exit
      -- CP-element group 381: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- CP-element group 381: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/$exit
      -- CP-element group 381: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_594/SplitProtocol/$exit
      -- CP-element group 381: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    phi_stmt_589_req_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_req_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(381), ack => phi_stmt_589_req_1); -- 
    checkNodeComputeEngine_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(379) & checkNodeComputeEngine_CP_1062_elements(380);
      gj_checkNodeComputeEngine_cp_element_group_381 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  transition  input  no-bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	376 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (2) 
      -- CP-element group 382: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Sample/ra
      -- 
    ra_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(382)); -- 
    -- CP-element group 383:  transition  input  no-bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	376 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (2) 
      -- CP-element group 383: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/Update/ca
      -- 
    ca_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (5) 
      -- CP-element group 384: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/$exit
      -- CP-element group 384: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$exit
      -- CP-element group 384: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/$exit
      -- CP-element group 384: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_604/SplitProtocol/$exit
      -- CP-element group 384: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_req
      -- 
    phi_stmt_599_req_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_599_req_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(384), ack => phi_stmt_599_req_1); -- 
    checkNodeComputeEngine_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(382) & checkNodeComputeEngine_CP_1062_elements(383);
      gj_checkNodeComputeEngine_cp_element_group_384 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  no-bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	378 
    -- CP-element group 385: 	381 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	406 
    -- CP-element group 385:  members (1) 
      -- CP-element group 385: 	 branch_block_stmt_226/bb_11_bb_14_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(378) & checkNodeComputeEngine_CP_1062_elements(381) & checkNodeComputeEngine_CP_1062_elements(384);
      gj_checkNodeComputeEngine_cp_element_group_385 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	213 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386: 	389 
    -- CP-element group 386: 	390 
    -- CP-element group 386: 	392 
    -- CP-element group 386: 	393 
    -- CP-element group 386:  members (19) 
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Sample/rr
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Update/cr
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Sample/rr
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Update/cr
      -- 
    rr_3199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(386), ack => type_cast_598_inst_req_0); -- 
    cr_3204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(386), ack => type_cast_598_inst_req_1); -- 
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(386), ack => type_cast_608_inst_req_0); -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(386), ack => type_cast_608_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(386) <= checkNodeComputeEngine_CP_1062_elements(213);
    -- CP-element group 387:  transition  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (1) 
      -- CP-element group 387: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_588_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(387) is a control-delay.
    cp_element_387_delay: control_delay_element  generic map(name => " 387_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(386), ack => checkNodeComputeEngine_CP_1062_elements(387), clk => clk, reset =>reset);
    -- CP-element group 388:  transition  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	395 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/$exit
      -- CP-element group 388: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$exit
      -- CP-element group 388: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_req
      -- 
    phi_stmt_576_req_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_576_req_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(388), ack => phi_stmt_576_req_3); -- 
    checkNodeComputeEngine_CP_1062_elements(388) <= checkNodeComputeEngine_CP_1062_elements(387);
    -- CP-element group 389:  transition  input  no-bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	386 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Sample/ra
      -- 
    ra_3200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(389)); -- 
    -- CP-element group 390:  transition  input  no-bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	386 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (2) 
      -- CP-element group 390: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/Update/ca
      -- 
    ca_3205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(390)); -- 
    -- CP-element group 391:  join  transition  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	395 
    -- CP-element group 391:  members (5) 
      -- CP-element group 391: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/$exit
      -- CP-element group 391: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- CP-element group 391: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/$exit
      -- CP-element group 391: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_598/SplitProtocol/$exit
      -- CP-element group 391: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    phi_stmt_589_req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(391), ack => phi_stmt_589_req_3); -- 
    checkNodeComputeEngine_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(389) & checkNodeComputeEngine_CP_1062_elements(390);
      gj_checkNodeComputeEngine_cp_element_group_391 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  transition  input  no-bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	386 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	394 
    -- CP-element group 392:  members (2) 
      -- CP-element group 392: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Sample/ra
      -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(392)); -- 
    -- CP-element group 393:  transition  input  no-bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	386 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (2) 
      -- CP-element group 393: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/Update/ca
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(393)); -- 
    -- CP-element group 394:  join  transition  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	392 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/$exit
      -- CP-element group 394: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$exit
      -- CP-element group 394: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/$exit
      -- CP-element group 394: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_608/SplitProtocol/$exit
      -- CP-element group 394: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_req
      -- 
    phi_stmt_599_req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_599_req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(394), ack => phi_stmt_599_req_3); -- 
    checkNodeComputeEngine_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(392) & checkNodeComputeEngine_CP_1062_elements(393);
      gj_checkNodeComputeEngine_cp_element_group_394 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  join  transition  no-bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	388 
    -- CP-element group 395: 	391 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	406 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 branch_block_stmt_226/bb_12_bb_14_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(388) & checkNodeComputeEngine_CP_1062_elements(391) & checkNodeComputeEngine_CP_1062_elements(394);
      gj_checkNodeComputeEngine_cp_element_group_395 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  fork  transition  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	26 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396: 	399 
    -- CP-element group 396: 	400 
    -- CP-element group 396: 	402 
    -- CP-element group 396: 	403 
    -- CP-element group 396:  members (19) 
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Update/cr
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Update/cr
      -- 
    rr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(396), ack => type_cast_596_inst_req_0); -- 
    cr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(396), ack => type_cast_596_inst_req_1); -- 
    rr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(396), ack => type_cast_606_inst_req_0); -- 
    cr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(396), ack => type_cast_606_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(396) <= checkNodeComputeEngine_CP_1062_elements(26);
    -- CP-element group 397:  transition  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/type_cast_585_konst_delay_trans
      -- 
    -- Element group checkNodeComputeEngine_CP_1062_elements(397) is a control-delay.
    cp_element_397_delay: control_delay_element  generic map(name => " 397_delay", delay_value => 1)  port map(req => checkNodeComputeEngine_CP_1062_elements(396), ack => checkNodeComputeEngine_CP_1062_elements(397), clk => clk, reset =>reset);
    -- CP-element group 398:  transition  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	405 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/$exit
      -- CP-element group 398: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_sources/$exit
      -- CP-element group 398: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_576/phi_stmt_576_req
      -- 
    phi_stmt_576_req_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_576_req_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(398), ack => phi_stmt_576_req_2); -- 
    checkNodeComputeEngine_CP_1062_elements(398) <= checkNodeComputeEngine_CP_1062_elements(397);
    -- CP-element group 399:  transition  input  no-bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	396 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	401 
    -- CP-element group 399:  members (2) 
      -- CP-element group 399: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Sample/ra
      -- 
    ra_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(399)); -- 
    -- CP-element group 400:  transition  input  no-bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	396 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/Update/ca
      -- 
    ca_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(400)); -- 
    -- CP-element group 401:  join  transition  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	399 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	405 
    -- CP-element group 401:  members (5) 
      -- CP-element group 401: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/$exit
      -- CP-element group 401: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- CP-element group 401: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/$exit
      -- CP-element group 401: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_596/SplitProtocol/$exit
      -- CP-element group 401: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    phi_stmt_589_req_3263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_req_3263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(401), ack => phi_stmt_589_req_2); -- 
    checkNodeComputeEngine_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(399) & checkNodeComputeEngine_CP_1062_elements(400);
      gj_checkNodeComputeEngine_cp_element_group_401 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  transition  input  no-bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	396 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (2) 
      -- CP-element group 402: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Sample/ra
      -- 
    ra_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(402)); -- 
    -- CP-element group 403:  transition  input  no-bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	396 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/Update/ca
      -- 
    ca_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(403)); -- 
    -- CP-element group 404:  join  transition  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (5) 
      -- CP-element group 404: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/$exit
      -- CP-element group 404: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/$exit
      -- CP-element group 404: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/$exit
      -- CP-element group 404: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_sources/type_cast_606/SplitProtocol/$exit
      -- CP-element group 404: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/phi_stmt_599/phi_stmt_599_req
      -- 
    phi_stmt_599_req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_599_req_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(404), ack => phi_stmt_599_req_2); -- 
    checkNodeComputeEngine_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(402) & checkNodeComputeEngine_CP_1062_elements(403);
      gj_checkNodeComputeEngine_cp_element_group_404 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  join  transition  no-bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	398 
    -- CP-element group 405: 	401 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (1) 
      -- CP-element group 405: 	 branch_block_stmt_226/bb_13_bb_14_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(398) & checkNodeComputeEngine_CP_1062_elements(401) & checkNodeComputeEngine_CP_1062_elements(404);
      gj_checkNodeComputeEngine_cp_element_group_405 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  merge  place  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	375 
    -- CP-element group 406: 	385 
    -- CP-element group 406: 	395 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (1) 
      -- CP-element group 406: 	 branch_block_stmt_226/merge_stmt_575_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(406) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(375) & checkNodeComputeEngine_CP_1062_elements(385) & checkNodeComputeEngine_CP_1062_elements(395) & checkNodeComputeEngine_CP_1062_elements(405));
    -- CP-element group 407:  fork  transition  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407: 	409 
    -- CP-element group 407: 	410 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_226/merge_stmt_575_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(407) <= checkNodeComputeEngine_CP_1062_elements(406);
    -- CP-element group 408:  transition  input  no-bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	411 
    -- CP-element group 408:  members (1) 
      -- CP-element group 408: 	 branch_block_stmt_226/merge_stmt_575_PhiAck/phi_stmt_576_ack
      -- 
    phi_stmt_576_ack_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_576_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(408)); -- 
    -- CP-element group 409:  transition  input  no-bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	407 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (1) 
      -- CP-element group 409: 	 branch_block_stmt_226/merge_stmt_575_PhiAck/phi_stmt_589_ack
      -- 
    phi_stmt_589_ack_3292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_589_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(409)); -- 
    -- CP-element group 410:  transition  input  no-bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	407 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (1) 
      -- CP-element group 410: 	 branch_block_stmt_226/merge_stmt_575_PhiAck/phi_stmt_599_ack
      -- 
    phi_stmt_599_ack_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_599_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(410)); -- 
    -- CP-element group 411:  join  transition  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	408 
    -- CP-element group 411: 	409 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	27 
    -- CP-element group 411:  members (1) 
      -- CP-element group 411: 	 branch_block_stmt_226/merge_stmt_575_PhiAck/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(408) & checkNodeComputeEngine_CP_1062_elements(409) & checkNodeComputeEngine_CP_1062_elements(410);
      gj_checkNodeComputeEngine_cp_element_group_411 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  fork  transition  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	226 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412: 	414 
    -- CP-element group 412: 	416 
    -- CP-element group 412: 	417 
    -- CP-element group 412:  members (17) 
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Sample/rr
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Update/cr
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Sample/rr
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Update/cr
      -- 
    rr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(412), ack => type_cast_631_inst_req_0); -- 
    cr_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(412), ack => type_cast_631_inst_req_1); -- 
    rr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(412), ack => type_cast_635_inst_req_0); -- 
    cr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(412), ack => type_cast_635_inst_req_1); -- 
    checkNodeComputeEngine_CP_1062_elements(412) <= checkNodeComputeEngine_CP_1062_elements(226);
    -- CP-element group 413:  transition  input  no-bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Sample/$exit
      -- CP-element group 413: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Sample/ra
      -- 
    ra_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(413)); -- 
    -- CP-element group 414:  transition  input  no-bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	412 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (2) 
      -- CP-element group 414: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/Update/ca
      -- 
    ca_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	413 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	419 
    -- CP-element group 415:  members (5) 
      -- CP-element group 415: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/$exit
      -- CP-element group 415: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/$exit
      -- CP-element group 415: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/$exit
      -- CP-element group 415: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_sources/type_cast_631/SplitProtocol/$exit
      -- CP-element group 415: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_628/phi_stmt_628_req
      -- 
    phi_stmt_628_req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_628_req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(415), ack => phi_stmt_628_req_0); -- 
    checkNodeComputeEngine_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(413) & checkNodeComputeEngine_CP_1062_elements(414);
      gj_checkNodeComputeEngine_cp_element_group_415 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  no-bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	412 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (2) 
      -- CP-element group 416: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Sample/ra
      -- 
    ra_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(416)); -- 
    -- CP-element group 417:  transition  input  no-bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	412 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (2) 
      -- CP-element group 417: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/Update/ca
      -- 
    ca_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_1, ack => checkNodeComputeEngine_CP_1062_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/$exit
      -- CP-element group 418: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/$exit
      -- CP-element group 418: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/$exit
      -- CP-element group 418: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_sources/type_cast_635/SplitProtocol/$exit
      -- CP-element group 418: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/phi_stmt_632/phi_stmt_632_req
      -- 
    phi_stmt_632_req_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_632_req_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => checkNodeComputeEngine_CP_1062_elements(418), ack => phi_stmt_632_req_0); -- 
    checkNodeComputeEngine_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(416) & checkNodeComputeEngine_CP_1062_elements(417);
      gj_checkNodeComputeEngine_cp_element_group_418 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  join  transition  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	415 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (1) 
      -- CP-element group 419: 	 branch_block_stmt_226/bb_14_xx_x_crit_edge_PhiReq/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(415) & checkNodeComputeEngine_CP_1062_elements(418);
      gj_checkNodeComputeEngine_cp_element_group_419 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  place  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (1) 
      -- CP-element group 420: 	 branch_block_stmt_226/merge_stmt_627_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(420) <= checkNodeComputeEngine_CP_1062_elements(419);
    -- CP-element group 421:  fork  transition  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421: 	423 
    -- CP-element group 421:  members (1) 
      -- CP-element group 421: 	 branch_block_stmt_226/merge_stmt_627_PhiAck/$entry
      -- 
    checkNodeComputeEngine_CP_1062_elements(421) <= checkNodeComputeEngine_CP_1062_elements(420);
    -- CP-element group 422:  transition  input  no-bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (1) 
      -- CP-element group 422: 	 branch_block_stmt_226/merge_stmt_627_PhiAck/phi_stmt_628_ack
      -- 
    phi_stmt_628_ack_3351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_628_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(422)); -- 
    -- CP-element group 423:  transition  input  no-bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (1) 
      -- CP-element group 423: 	 branch_block_stmt_226/merge_stmt_627_PhiAck/phi_stmt_632_ack
      -- 
    phi_stmt_632_ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_632_ack_0, ack => checkNodeComputeEngine_CP_1062_elements(423)); -- 
    -- CP-element group 424:  join  transition  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	29 
    -- CP-element group 424:  members (1) 
      -- CP-element group 424: 	 branch_block_stmt_226/merge_stmt_627_PhiAck/$exit
      -- 
    checkNodeComputeEngine_cp_element_group_424: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "checkNodeComputeEngine_cp_element_group_424"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= checkNodeComputeEngine_CP_1062_elements(422) & checkNodeComputeEngine_CP_1062_elements(423);
      gj_checkNodeComputeEngine_cp_element_group_424 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => checkNodeComputeEngine_CP_1062_elements(424), clk => clk, reset => reset); --
    end block;
    -- CP-element group 425:  transition  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	254 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (2) 
      -- CP-element group 425: 	 branch_block_stmt_226/xx_x_crit_edge_xx_x_crit_edge9x_xloopexit_PhiReq/$entry
      -- CP-element group 425: 	 branch_block_stmt_226/xx_x_crit_edge_xx_x_crit_edge9x_xloopexit_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(425) <= checkNodeComputeEngine_CP_1062_elements(254);
    -- CP-element group 426:  place  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (1) 
      -- CP-element group 426: 	 branch_block_stmt_226/merge_stmt_686_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(426) <= checkNodeComputeEngine_CP_1062_elements(425);
    -- CP-element group 427:  transition  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	31 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_226/merge_stmt_686_PhiAck/$entry
      -- CP-element group 427: 	 branch_block_stmt_226/merge_stmt_686_PhiAck/$exit
      -- CP-element group 427: 	 branch_block_stmt_226/merge_stmt_686_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(427) <= checkNodeComputeEngine_CP_1062_elements(426);
    -- CP-element group 428:  transition  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	126 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	430 
    -- CP-element group 428:  members (2) 
      -- CP-element group 428: 	 branch_block_stmt_226/bb_5_xx_x_crit_edge9_PhiReq/$entry
      -- CP-element group 428: 	 branch_block_stmt_226/bb_5_xx_x_crit_edge9_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(428) <= checkNodeComputeEngine_CP_1062_elements(126);
    -- CP-element group 429:  transition  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	31 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (2) 
      -- CP-element group 429: 	 branch_block_stmt_226/xx_x_crit_edge9x_xloopexit_xx_x_crit_edge9_PhiReq/$entry
      -- CP-element group 429: 	 branch_block_stmt_226/xx_x_crit_edge9x_xloopexit_xx_x_crit_edge9_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(429) <= checkNodeComputeEngine_CP_1062_elements(31);
    -- CP-element group 430:  merge  place  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	428 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (1) 
      -- CP-element group 430: 	 branch_block_stmt_226/merge_stmt_688_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(430) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(428) & checkNodeComputeEngine_CP_1062_elements(429));
    -- CP-element group 431:  transition  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	32 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_226/merge_stmt_688_PhiAck/$entry
      -- CP-element group 431: 	 branch_block_stmt_226/merge_stmt_688_PhiAck/$exit
      -- CP-element group 431: 	 branch_block_stmt_226/merge_stmt_688_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(431) <= checkNodeComputeEngine_CP_1062_elements(430);
    -- CP-element group 432:  transition  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	267 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (2) 
      -- CP-element group 432: 	 branch_block_stmt_226/xx_x_crit_edge9_xx_x_crit_edge12x_xloopexit_PhiReq/$entry
      -- CP-element group 432: 	 branch_block_stmt_226/xx_x_crit_edge9_xx_x_crit_edge12x_xloopexit_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(432) <= checkNodeComputeEngine_CP_1062_elements(267);
    -- CP-element group 433:  place  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (1) 
      -- CP-element group 433: 	 branch_block_stmt_226/merge_stmt_700_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(433) <= checkNodeComputeEngine_CP_1062_elements(432);
    -- CP-element group 434:  transition  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	34 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_226/merge_stmt_700_PhiAck/$entry
      -- CP-element group 434: 	 branch_block_stmt_226/merge_stmt_700_PhiAck/$exit
      -- CP-element group 434: 	 branch_block_stmt_226/merge_stmt_700_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(434) <= checkNodeComputeEngine_CP_1062_elements(433);
    -- CP-element group 435:  transition  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	49 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	437 
    -- CP-element group 435:  members (2) 
      -- CP-element group 435: 	 branch_block_stmt_226/bb_0_xx_x_crit_edge12_PhiReq/$entry
      -- CP-element group 435: 	 branch_block_stmt_226/bb_0_xx_x_crit_edge12_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(435) <= checkNodeComputeEngine_CP_1062_elements(49);
    -- CP-element group 436:  transition  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	34 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (2) 
      -- CP-element group 436: 	 branch_block_stmt_226/xx_x_crit_edge12x_xloopexit_xx_x_crit_edge12_PhiReq/$entry
      -- CP-element group 436: 	 branch_block_stmt_226/xx_x_crit_edge12x_xloopexit_xx_x_crit_edge12_PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(436) <= checkNodeComputeEngine_CP_1062_elements(34);
    -- CP-element group 437:  merge  place  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	435 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (1) 
      -- CP-element group 437: 	 branch_block_stmt_226/merge_stmt_702_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(437) <= OrReduce(checkNodeComputeEngine_CP_1062_elements(435) & checkNodeComputeEngine_CP_1062_elements(436));
    -- CP-element group 438:  transition  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	35 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_226/merge_stmt_702_PhiAck/$entry
      -- CP-element group 438: 	 branch_block_stmt_226/merge_stmt_702_PhiAck/$exit
      -- CP-element group 438: 	 branch_block_stmt_226/merge_stmt_702_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(438) <= checkNodeComputeEngine_CP_1062_elements(437);
    -- CP-element group 439:  transition  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	35 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (2) 
      -- CP-element group 439: 	 branch_block_stmt_226/return___PhiReq/$entry
      -- CP-element group 439: 	 branch_block_stmt_226/return___PhiReq/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(439) <= checkNodeComputeEngine_CP_1062_elements(35);
    -- CP-element group 440:  place  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (1) 
      -- CP-element group 440: 	 branch_block_stmt_226/merge_stmt_704_PhiReqMerge
      -- 
    checkNodeComputeEngine_CP_1062_elements(440) <= checkNodeComputeEngine_CP_1062_elements(439);
    -- CP-element group 441:  transition  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	36 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_226/merge_stmt_704_PhiAck/$entry
      -- CP-element group 441: 	 branch_block_stmt_226/merge_stmt_704_PhiAck/$exit
      -- CP-element group 441: 	 branch_block_stmt_226/merge_stmt_704_PhiAck/dummy
      -- 
    checkNodeComputeEngine_CP_1062_elements(441) <= checkNodeComputeEngine_CP_1062_elements(440);
    -- CP-element group 442:  transition  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	36 
    -- CP-element group 442: successors 
    -- CP-element group 442:  members (2) 
      -- CP-element group 442: 	 $exit
      -- CP-element group 442: 	 branch_block_stmt_226/$exit
      -- 
    checkNodeComputeEngine_CP_1062_elements(442) <= checkNodeComputeEngine_CP_1062_elements(36);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_ncol_ind_266_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncol_ind_266_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_nrows_228_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_nrows_228_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_nrows_274_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_nrows_274_word_address_0 : std_logic_vector(0 downto 0);
    signal R_iNsTr_17_329_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_17_329_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_17_354_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_17_354_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_24_334_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_24_334_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_37_411_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_37_411_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_45_482_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_45_482_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_63_661_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_63_661_scaled : std_logic_vector(9 downto 0);
    signal array_obj_ref_330_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_330_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_330_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_330_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_335_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_335_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_335_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_335_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_355_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_355_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_355_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_355_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_412_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_412_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_412_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_412_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_483_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_483_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_483_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_483_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_662_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_662_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_662_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_662_root_address : std_logic_vector(9 downto 0);
    signal exitcond1_620 : std_logic_vector(0 downto 0);
    signal exitcond_679 : std_logic_vector(0 downto 0);
    signal exorx_x0_548 : std_logic_vector(7 downto 0);
    signal exorx_x1_599 : std_logic_vector(7 downto 0);
    signal exorx_x1x_xlcssa_628 : std_logic_vector(7 downto 0);
    signal exorx_x25_442 : std_logic_vector(7 downto 0);
    signal flagx_x0_576 : std_logic_vector(7 downto 0);
    signal flagx_x12_464 : std_logic_vector(7 downto 0);
    signal iNsTr_0_229 : std_logic_vector(15 downto 0);
    signal iNsTr_10_275 : std_logic_vector(15 downto 0);
    signal iNsTr_11_279 : std_logic_vector(31 downto 0);
    signal iNsTr_12_285 : std_logic_vector(31 downto 0);
    signal iNsTr_13_290 : std_logic_vector(0 downto 0);
    signal iNsTr_14_294 : std_logic_vector(63 downto 0);
    signal iNsTr_15_298 : std_logic_vector(63 downto 0);
    signal iNsTr_16_304 : std_logic_vector(63 downto 0);
    signal iNsTr_17_309 : std_logic_vector(63 downto 0);
    signal iNsTr_19_357 : std_logic_vector(31 downto 0);
    signal iNsTr_1_235 : std_logic_vector(0 downto 0);
    signal iNsTr_20_361 : std_logic_vector(15 downto 0);
    signal iNsTr_21_372 : std_logic_vector(15 downto 0);
    signal iNsTr_23_322 : std_logic_vector(63 downto 0);
    signal iNsTr_24_327 : std_logic_vector(63 downto 0);
    signal iNsTr_25_332 : std_logic_vector(31 downto 0);
    signal iNsTr_26_337 : std_logic_vector(31 downto 0);
    signal iNsTr_27_341 : std_logic_vector(15 downto 0);
    signal iNsTr_28_345 : std_logic_vector(15 downto 0);
    signal iNsTr_29_350 : std_logic_vector(15 downto 0);
    signal iNsTr_31_387 : std_logic_vector(0 downto 0);
    signal iNsTr_33_693 : std_logic_vector(0 downto 0);
    signal iNsTr_35_398 : std_logic_vector(63 downto 0);
    signal iNsTr_36_404 : std_logic_vector(63 downto 0);
    signal iNsTr_37_409 : std_logic_vector(63 downto 0);
    signal iNsTr_38_414 : std_logic_vector(31 downto 0);
    signal iNsTr_39_418 : std_logic_vector(15 downto 0);
    signal iNsTr_42_427 : std_logic_vector(15 downto 0);
    signal iNsTr_44_450 : std_logic_vector(15 downto 0);
    signal iNsTr_45_480 : std_logic_vector(63 downto 0);
    signal iNsTr_46_485 : std_logic_vector(31 downto 0);
    signal iNsTr_47_489 : std_logic_vector(31 downto 0);
    signal iNsTr_48_493 : std_logic_vector(63 downto 0);
    signal iNsTr_49_499 : std_logic_vector(0 downto 0);
    signal iNsTr_51_512 : std_logic_vector(31 downto 0);
    signal iNsTr_53_526 : std_logic_vector(0 downto 0);
    signal iNsTr_55_615 : std_logic_vector(15 downto 0);
    signal iNsTr_57_539 : std_logic_vector(0 downto 0);
    signal iNsTr_58_543 : std_logic_vector(7 downto 0);
    signal iNsTr_59_554 : std_logic_vector(0 downto 0);
    signal iNsTr_5_245 : std_logic_vector(15 downto 0);
    signal iNsTr_61_642 : std_logic_vector(0 downto 0);
    signal iNsTr_62_655 : std_logic_vector(31 downto 0);
    signal iNsTr_63_659 : std_logic_vector(63 downto 0);
    signal iNsTr_64_664 : std_logic_vector(31 downto 0);
    signal iNsTr_66_674 : std_logic_vector(15 downto 0);
    signal iNsTr_68_566 : std_logic_vector(0 downto 0);
    signal iNsTr_6_264 : std_logic_vector(15 downto 0);
    signal iNsTr_8_267 : std_logic_vector(15 downto 0);
    signal iNsTr_9_272 : std_logic_vector(31 downto 0);
    signal ptr_deref_340_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_340_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_340_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_340_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_340_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_344_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_344_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_344_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_344_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_344_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_360_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_360_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_360_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_360_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_360_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_417_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_417_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_417_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_417_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_417_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_488_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_488_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_488_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_488_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_488_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_666_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_666_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_666_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_666_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_666_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_666_word_offset_0 : std_logic_vector(9 downto 0);
    signal rangex_x0_375 : std_logic_vector(15 downto 0);
    signal signx_x0_650 : std_logic_vector(31 downto 0);
    signal temp1x_x0_515 : std_logic_vector(31 downto 0);
    signal tmp13_476 : std_logic_vector(15 downto 0);
    signal tmp15_424 : std_logic_vector(15 downto 0);
    signal tmp16_439 : std_logic_vector(15 downto 0);
    signal tmp17_258 : std_logic_vector(15 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_248_wire : std_logic_vector(15 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_256_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_262_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_283_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_302_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_365_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_378_wire : std_logic_vector(15 downto 0);
    signal type_cast_380_wire : std_logic_vector(15 downto 0);
    signal type_cast_385_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_402_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_422_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_431_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_433_wire : std_logic_vector(15 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_449_wire : std_logic_vector(7 downto 0);
    signal type_cast_454_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_456_wire : std_logic_vector(15 downto 0);
    signal type_cast_461_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_463_wire : std_logic_vector(31 downto 0);
    signal type_cast_468_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_470_wire : std_logic_vector(7 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_509_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_518_wire : std_logic_vector(31 downto 0);
    signal type_cast_520_wire : std_logic_vector(31 downto 0);
    signal type_cast_537_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_552_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_579_wire : std_logic_vector(7 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_585_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_592_wire : std_logic_vector(31 downto 0);
    signal type_cast_594_wire : std_logic_vector(31 downto 0);
    signal type_cast_596_wire : std_logic_vector(31 downto 0);
    signal type_cast_598_wire : std_logic_vector(31 downto 0);
    signal type_cast_602_wire : std_logic_vector(7 downto 0);
    signal type_cast_604_wire : std_logic_vector(7 downto 0);
    signal type_cast_606_wire : std_logic_vector(7 downto 0);
    signal type_cast_608_wire : std_logic_vector(7 downto 0);
    signal type_cast_613_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_631_wire : std_logic_vector(7 downto 0);
    signal type_cast_635_wire : std_logic_vector(31 downto 0);
    signal type_cast_640_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_646_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_672_wire_constant : std_logic_vector(15 downto 0);
    signal valx_x1_589 : std_logic_vector(31 downto 0);
    signal valx_x1x_xlcssa_632 : std_logic_vector(31 downto 0);
    signal valx_x23_457 : std_logic_vector(31 downto 0);
    signal xx_xneg1_367 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_ncol_ind_266_word_address_0 <= "0";
    LOAD_nrows_228_word_address_0 <= "0";
    LOAD_nrows_274_word_address_0 <= "0";
    array_obj_ref_330_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_330_resized_base_address <= "0000000000";
    array_obj_ref_335_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_335_resized_base_address <= "0000000000";
    array_obj_ref_355_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_355_resized_base_address <= "0000000000";
    array_obj_ref_412_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_412_resized_base_address <= "0000000000";
    array_obj_ref_483_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_483_resized_base_address <= "0000000000";
    array_obj_ref_662_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_662_resized_base_address <= "0000000000";
    ptr_deref_340_word_offset_0 <= "0000000000";
    ptr_deref_344_word_offset_0 <= "0000000000";
    ptr_deref_360_word_offset_0 <= "0000000000";
    ptr_deref_417_word_offset_0 <= "0000000000";
    ptr_deref_488_word_offset_0 <= "0000000000";
    ptr_deref_666_word_offset_0 <= "0000000000";
    type_cast_233_wire_constant <= "0000000000000000";
    type_cast_251_wire_constant <= "0000000000000000";
    type_cast_256_wire_constant <= "0000000000000001";
    type_cast_262_wire_constant <= "0000000000000001";
    type_cast_283_wire_constant <= "11111111111111111111111111111111";
    type_cast_302_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_320_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_365_wire_constant <= "0000000000000001";
    type_cast_385_wire_constant <= "0000000000000000";
    type_cast_402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_422_wire_constant <= "1111111111111111";
    type_cast_431_wire_constant <= "0000000000000000";
    type_cast_447_wire_constant <= "00000000";
    type_cast_454_wire_constant <= "0000000000000000";
    type_cast_461_wire_constant <= "00000000000000000000000000000000";
    type_cast_468_wire_constant <= "00000000";
    type_cast_497_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_509_wire_constant <= "10000000000000000000000000000000";
    type_cast_537_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_552_wire_constant <= "00000000";
    type_cast_582_wire_constant <= "00000001";
    type_cast_585_wire_constant <= "00000001";
    type_cast_588_wire_constant <= "00000001";
    type_cast_613_wire_constant <= "0000000000000001";
    type_cast_640_wire_constant <= "00000000";
    type_cast_646_wire_constant <= "00111111100000000000000000000000";
    type_cast_648_wire_constant <= "10111111100000000000000000000000";
    type_cast_672_wire_constant <= "0000000000000001";
    phi_stmt_245: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_248_wire & type_cast_251_wire_constant;
      req <= phi_stmt_245_req_0 & phi_stmt_245_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_245",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_245_ack_0,
          idata => idata,
          odata => iNsTr_5_245,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_245
    phi_stmt_375: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_378_wire & type_cast_380_wire;
      req <= phi_stmt_375_req_0 & phi_stmt_375_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_375",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_375_ack_0,
          idata => idata,
          odata => rangex_x0_375,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_375
    phi_stmt_427: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_431_wire_constant & type_cast_433_wire;
      req <= phi_stmt_427_req_0 & phi_stmt_427_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_427",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_427_ack_0,
          idata => idata,
          odata => iNsTr_42_427,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_427
    phi_stmt_442: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_447_wire_constant & type_cast_449_wire;
      req <= phi_stmt_442_req_0 & phi_stmt_442_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_442",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_442_ack_0,
          idata => idata,
          odata => exorx_x25_442,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_442
    phi_stmt_450: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_454_wire_constant & type_cast_456_wire;
      req <= phi_stmt_450_req_0 & phi_stmt_450_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_450",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_450_ack_0,
          idata => idata,
          odata => iNsTr_44_450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_450
    phi_stmt_457: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_461_wire_constant & type_cast_463_wire;
      req <= phi_stmt_457_req_0 & phi_stmt_457_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_457",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_457_ack_0,
          idata => idata,
          odata => valx_x23_457,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_457
    phi_stmt_464: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_468_wire_constant & type_cast_470_wire;
      req <= phi_stmt_464_req_0 & phi_stmt_464_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_464",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_464_ack_0,
          idata => idata,
          odata => flagx_x12_464,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_464
    phi_stmt_515: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_518_wire & type_cast_520_wire;
      req <= phi_stmt_515_req_0 & phi_stmt_515_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_515",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_515_ack_0,
          idata => idata,
          odata => temp1x_x0_515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_515
    phi_stmt_576: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(3 downto 0);
      --
    begin -- 
      idata <= type_cast_579_wire & type_cast_582_wire_constant & type_cast_585_wire_constant & type_cast_588_wire_constant;
      req <= phi_stmt_576_req_0 & phi_stmt_576_req_1 & phi_stmt_576_req_2 & phi_stmt_576_req_3;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_576",
          num_reqs => 4,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_576_ack_0,
          idata => idata,
          odata => flagx_x0_576,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_576
    phi_stmt_589: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(3 downto 0);
      --
    begin -- 
      idata <= type_cast_592_wire & type_cast_594_wire & type_cast_596_wire & type_cast_598_wire;
      req <= phi_stmt_589_req_0 & phi_stmt_589_req_1 & phi_stmt_589_req_2 & phi_stmt_589_req_3;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_589",
          num_reqs => 4,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_589_ack_0,
          idata => idata,
          odata => valx_x1_589,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_589
    phi_stmt_599: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(3 downto 0);
      --
    begin -- 
      idata <= type_cast_602_wire & type_cast_604_wire & type_cast_606_wire & type_cast_608_wire;
      req <= phi_stmt_599_req_0 & phi_stmt_599_req_1 & phi_stmt_599_req_2 & phi_stmt_599_req_3;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_599",
          num_reqs => 4,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_599_ack_0,
          idata => idata,
          odata => exorx_x1_599,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_599
    phi_stmt_628: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_631_wire;
      req(0) <= phi_stmt_628_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_628",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_628_ack_0,
          idata => idata,
          odata => exorx_x1x_xlcssa_628,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_628
    phi_stmt_632: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_635_wire;
      req(0) <= phi_stmt_632_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_632",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_632_ack_0,
          idata => idata,
          odata => valx_x1x_xlcssa_632,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_632
    MUX_649_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_649_inst_req_0;
      MUX_649_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_649_inst_req_1;
      MUX_649_inst_ack_1<= update_ack(0);
      MUX_649_inst: SelectSplitProtocol generic map(name => "MUX_649_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_646_wire_constant, y => type_cast_648_wire_constant, sel => iNsTr_61_642, z => signx_x0_650, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    addr_of_331_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_331_final_reg_req_0;
      addr_of_331_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_331_final_reg_req_1;
      addr_of_331_final_reg_ack_1<= rack(0);
      addr_of_331_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_331_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_330_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_25_332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_336_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_336_final_reg_req_0;
      addr_of_336_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_336_final_reg_req_1;
      addr_of_336_final_reg_ack_1<= rack(0);
      addr_of_336_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_336_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_335_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_356_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_356_final_reg_req_0;
      addr_of_356_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_356_final_reg_req_1;
      addr_of_356_final_reg_ack_1<= rack(0);
      addr_of_356_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_356_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_355_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_413_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_413_final_reg_req_0;
      addr_of_413_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_413_final_reg_req_1;
      addr_of_413_final_reg_ack_1<= rack(0);
      addr_of_413_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_413_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_412_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_38_414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_484_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_484_final_reg_req_0;
      addr_of_484_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_484_final_reg_req_1;
      addr_of_484_final_reg_ack_1<= rack(0);
      addr_of_484_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_484_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_483_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_46_485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_663_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_663_final_reg_req_0;
      addr_of_663_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_663_final_reg_req_1;
      addr_of_663_final_reg_ack_1<= rack(0);
      addr_of_663_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_663_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_662_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_64_664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_248_inst_req_0;
      type_cast_248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_248_inst_req_1;
      type_cast_248_inst_ack_1<= rack(0);
      type_cast_248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_6_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_248_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_271_inst_req_0;
      type_cast_271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_271_inst_req_1;
      type_cast_271_inst_ack_1<= rack(0);
      type_cast_271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_5_245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_9_272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_278_inst_req_0;
      type_cast_278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_278_inst_req_1;
      type_cast_278_inst_ack_1<= rack(0);
      type_cast_278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_10_275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_11_279,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_293_inst_req_0;
      type_cast_293_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_293_inst_req_1;
      type_cast_293_inst_ack_1<= rack(0);
      type_cast_293_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_293_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_8_267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_294,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_297_inst_req_0;
      type_cast_297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_297_inst_req_1;
      type_cast_297_inst_ack_1<= rack(0);
      type_cast_297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_5_245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_15_298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_378_inst_req_0;
      type_cast_378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_378_inst_req_1;
      type_cast_378_inst_ack_1<= rack(0);
      type_cast_378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_21_372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_378_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_29_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_380_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_397_inst_req_0;
      type_cast_397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_397_inst_req_1;
      type_cast_397_inst_ack_1<= rack(0);
      type_cast_397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_5_245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_35_398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_433_inst_req_0;
      type_cast_433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_433_inst_req_1;
      type_cast_433_inst_ack_1<= rack(0);
      type_cast_433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_66_674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_433_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_449_inst_req_0;
      type_cast_449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_449_inst_req_1;
      type_cast_449_inst_ack_1<= rack(0);
      type_cast_449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x1_599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_449_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_55_615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_456_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_463_inst_req_0;
      type_cast_463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_463_inst_req_1;
      type_cast_463_inst_ack_1<= rack(0);
      type_cast_463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valx_x1_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_463_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_470_inst_req_0;
      type_cast_470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_470_inst_req_1;
      type_cast_470_inst_ack_1<= rack(0);
      type_cast_470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => flagx_x0_576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_470_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_479_inst_req_0;
      type_cast_479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_479_inst_req_1;
      type_cast_479_inst_ack_1<= rack(0);
      type_cast_479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp13_476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_45_480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_518_inst_req_0;
      type_cast_518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_518_inst_req_1;
      type_cast_518_inst_ack_1<= rack(0);
      type_cast_518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_51_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_518_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_47_489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_520_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_542_inst_req_0;
      type_cast_542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_542_inst_req_1;
      type_cast_542_inst_ack_1<= rack(0);
      type_cast_542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_57_539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_58_543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_579_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_579_inst_req_0;
      type_cast_579_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_579_inst_req_1;
      type_cast_579_inst_ack_1<= rack(0);
      type_cast_579_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_579_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => flagx_x12_464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_579_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valx_x23_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_592_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_594_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_594_inst_req_0;
      type_cast_594_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_594_inst_req_1;
      type_cast_594_inst_ack_1<= rack(0);
      type_cast_594_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_594_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => temp1x_x0_515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_594_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_596_inst_req_0;
      type_cast_596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_596_inst_req_1;
      type_cast_596_inst_ack_1<= rack(0);
      type_cast_596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => temp1x_x0_515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_596_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valx_x23_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_598_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_602_inst_req_0;
      type_cast_602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_602_inst_req_1;
      type_cast_602_inst_ack_1<= rack(0);
      type_cast_602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x25_442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_602_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_604_inst_req_0;
      type_cast_604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_604_inst_req_1;
      type_cast_604_inst_ack_1<= rack(0);
      type_cast_604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x0_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_604_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_606_inst_req_0;
      type_cast_606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_606_inst_req_1;
      type_cast_606_inst_ack_1<= rack(0);
      type_cast_606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x0_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x0_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_608_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exorx_x1_599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_631_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_635_inst_req_0;
      type_cast_635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_635_inst_req_1;
      type_cast_635_inst_ack_1<= rack(0);
      type_cast_635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valx_x1_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_635_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_658_inst_req_0;
      type_cast_658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_658_inst_req_1;
      type_cast_658_inst_ack_1<= rack(0);
      type_cast_658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_63_659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_ncol_ind_266_gather_scatter
    process(LOAD_ncol_ind_266_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncol_ind_266_data_0;
      ov(15 downto 0) := iv;
      iNsTr_8_267 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_nrows_228_gather_scatter
    process(LOAD_nrows_228_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_nrows_228_data_0;
      ov(15 downto 0) := iv;
      iNsTr_0_229 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_nrows_274_gather_scatter
    process(LOAD_nrows_274_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_nrows_274_data_0;
      ov(15 downto 0) := iv;
      iNsTr_10_275 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_330_index_0_rename
    process(R_iNsTr_17_329_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_17_329_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_17_329_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_330_index_0_resize
    process(iNsTr_17_309) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_309;
      ov := iv(9 downto 0);
      R_iNsTr_17_329_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_330_index_offset
    process(R_iNsTr_17_329_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_17_329_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_330_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_330_root_address_inst
    process(array_obj_ref_330_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_330_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_330_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_index_0_rename
    process(R_iNsTr_24_334_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_24_334_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_24_334_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_index_0_resize
    process(iNsTr_24_327) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_24_327;
      ov := iv(9 downto 0);
      R_iNsTr_24_334_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_index_offset
    process(R_iNsTr_24_334_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_24_334_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_335_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_root_address_inst
    process(array_obj_ref_335_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_335_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_335_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_index_0_rename
    process(R_iNsTr_17_354_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_17_354_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_17_354_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_index_0_resize
    process(iNsTr_17_309) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_309;
      ov := iv(9 downto 0);
      R_iNsTr_17_354_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_index_offset
    process(R_iNsTr_17_354_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_17_354_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_355_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_root_address_inst
    process(array_obj_ref_355_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_355_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_355_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_index_0_rename
    process(R_iNsTr_37_411_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_37_411_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_37_411_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_index_0_resize
    process(iNsTr_37_409) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_409;
      ov := iv(9 downto 0);
      R_iNsTr_37_411_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_index_offset
    process(R_iNsTr_37_411_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_37_411_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_412_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_root_address_inst
    process(array_obj_ref_412_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_412_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_412_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_index_0_rename
    process(R_iNsTr_45_482_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_45_482_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_45_482_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_index_0_resize
    process(iNsTr_45_480) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_45_480;
      ov := iv(9 downto 0);
      R_iNsTr_45_482_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_index_offset
    process(R_iNsTr_45_482_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_45_482_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_483_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_483_root_address_inst
    process(array_obj_ref_483_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_483_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_483_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_662_index_0_rename
    process(R_iNsTr_63_661_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_63_661_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_63_661_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_662_index_0_resize
    process(iNsTr_63_659) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_63_659;
      ov := iv(9 downto 0);
      R_iNsTr_63_661_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_662_index_offset
    process(R_iNsTr_63_661_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_63_661_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_662_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_662_root_address_inst
    process(array_obj_ref_662_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_662_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_662_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_addr_0
    process(ptr_deref_340_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_340_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_base_resize
    process(iNsTr_25_332) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_332;
      ov := iv(9 downto 0);
      ptr_deref_340_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_gather_scatter
    process(ptr_deref_340_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_data_0;
      ov(15 downto 0) := iv;
      iNsTr_27_341 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_root_address_inst
    process(ptr_deref_340_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_340_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_344_addr_0
    process(ptr_deref_344_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_344_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_344_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_344_base_resize
    process(iNsTr_26_337) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_337;
      ov := iv(9 downto 0);
      ptr_deref_344_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_344_gather_scatter
    process(ptr_deref_344_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_344_data_0;
      ov(15 downto 0) := iv;
      iNsTr_28_345 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_344_root_address_inst
    process(ptr_deref_344_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_344_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_344_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_360_addr_0
    process(ptr_deref_360_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_360_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_360_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_360_base_resize
    process(iNsTr_19_357) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_357;
      ov := iv(9 downto 0);
      ptr_deref_360_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_360_gather_scatter
    process(ptr_deref_360_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_360_data_0;
      ov(15 downto 0) := iv;
      iNsTr_20_361 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_360_root_address_inst
    process(ptr_deref_360_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_360_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_360_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_417_addr_0
    process(ptr_deref_417_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_417_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_417_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_417_base_resize
    process(iNsTr_38_414) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_414;
      ov := iv(9 downto 0);
      ptr_deref_417_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_417_gather_scatter
    process(ptr_deref_417_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_417_data_0;
      ov(15 downto 0) := iv;
      iNsTr_39_418 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_417_root_address_inst
    process(ptr_deref_417_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_417_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_417_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_addr_0
    process(ptr_deref_488_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_488_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_base_resize
    process(iNsTr_46_485) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_485;
      ov := iv(9 downto 0);
      ptr_deref_488_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_gather_scatter
    process(ptr_deref_488_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_data_0;
      ov(31 downto 0) := iv;
      iNsTr_47_489 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_488_root_address_inst
    process(ptr_deref_488_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_488_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_488_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_addr_0
    process(ptr_deref_666_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_666_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_666_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_base_resize
    process(iNsTr_64_664) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_64_664;
      ov := iv(9 downto 0);
      ptr_deref_666_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_gather_scatter
    process(iNsTr_62_655) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_62_655;
      ov(31 downto 0) := iv;
      ptr_deref_666_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_666_root_address_inst
    process(ptr_deref_666_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_666_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_666_root_address <= ov(9 downto 0);
      --
    end process;
    if_stmt_236_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_1_235;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_236_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_236_branch_req_0,
          ack0 => if_stmt_236_branch_ack_0,
          ack1 => if_stmt_236_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_310_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_13_290;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_310_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_310_branch_req_0,
          ack0 => if_stmt_310_branch_ack_0,
          ack1 => if_stmt_310_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_388_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_31_387;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_388_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_388_branch_req_0,
          ack0 => if_stmt_388_branch_ack_0,
          ack1 => if_stmt_388_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_500_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_49_499;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_500_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_500_branch_req_0,
          ack0 => if_stmt_500_branch_ack_0,
          ack1 => if_stmt_500_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_527_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_53_526;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_527_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_527_branch_req_0,
          ack0 => if_stmt_527_branch_ack_0,
          ack1 => if_stmt_527_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_555_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_59_554;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_555_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_555_branch_req_0,
          ack0 => if_stmt_555_branch_ack_0,
          ack1 => if_stmt_555_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_567_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_68_566;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_567_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_567_branch_req_0,
          ack0 => if_stmt_567_branch_ack_0,
          ack1 => if_stmt_567_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_621_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_620;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_621_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_621_branch_req_0,
          ack0 => if_stmt_621_branch_ack_0,
          ack1 => if_stmt_621_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_680_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_679;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_680_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_680_branch_req_0,
          ack0 => if_stmt_680_branch_ack_0,
          ack1 => if_stmt_680_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_694_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_33_693;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_694_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_694_branch_req_0,
          ack0 => if_stmt_694_branch_ack_0,
          ack1 => if_stmt_694_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u16_u16_257_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_5_245;
      tmp17_258 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_257_inst_req_0;
      ADD_u16_u16_257_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_257_inst_req_1;
      ADD_u16_u16_257_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u16_u16_263_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_5_245;
      iNsTr_6_264 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_263_inst_req_0;
      ADD_u16_u16_263_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_263_inst_req_1;
      ADD_u16_u16_263_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u16_u16_366_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_8_267;
      xx_xneg1_367 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_366_inst_req_0;
      ADD_u16_u16_366_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_366_inst_req_1;
      ADD_u16_u16_366_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u16_u16_423_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_39_418;
      tmp15_424 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_423_inst_req_0;
      ADD_u16_u16_423_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_423_inst_req_1;
      ADD_u16_u16_423_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ADD_u16_u16_438_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp15_424 & iNsTr_42_427;
      tmp16_439 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_438_inst_req_0;
      ADD_u16_u16_438_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_438_inst_req_1;
      ADD_u16_u16_438_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ADD_u16_u16_475_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp15_424 & iNsTr_44_450;
      tmp13_476 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_475_inst_req_0;
      ADD_u16_u16_475_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_475_inst_req_1;
      ADD_u16_u16_475_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : ADD_u16_u16_614_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_44_450;
      iNsTr_55_615 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_614_inst_req_0;
      ADD_u16_u16_614_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_614_inst_req_1;
      ADD_u16_u16_614_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ADD_u16_u16_673_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_42_427;
      iNsTr_66_674 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_673_inst_req_0;
      ADD_u16_u16_673_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_673_inst_req_1;
      ADD_u16_u16_673_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ADD_u32_u32_284_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_11_279;
      iNsTr_12_285 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_284_inst_req_0;
      ADD_u32_u32_284_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_284_inst_req_1;
      ADD_u32_u32_284_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_8_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ADD_u64_u64_303_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_15_298;
      iNsTr_16_304 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_303_inst_req_0;
      ADD_u64_u64_303_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_303_inst_req_1;
      ADD_u64_u64_303_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_9_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ADD_u64_u64_308_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_16_304 & iNsTr_14_294;
      iNsTr_17_309 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_308_inst_req_0;
      ADD_u64_u64_308_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_308_inst_req_1;
      ADD_u64_u64_308_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_10_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ADD_u64_u64_321_inst 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_15_298;
      iNsTr_23_322 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_321_inst_req_0;
      ADD_u64_u64_321_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_321_inst_req_1;
      ADD_u64_u64_321_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000100",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ADD_u64_u64_326_inst 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_23_322 & iNsTr_14_294;
      iNsTr_24_327 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_326_inst_req_0;
      ADD_u64_u64_326_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_326_inst_req_1;
      ADD_u64_u64_326_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_12_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ADD_u64_u64_403_inst 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_35_398;
      iNsTr_36_404 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_403_inst_req_0;
      ADD_u64_u64_403_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_403_inst_req_1;
      ADD_u64_u64_403_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ADD_u64_u64_408_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_36_404 & iNsTr_14_294;
      iNsTr_37_409 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_408_inst_req_0;
      ADD_u64_u64_408_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_408_inst_req_1;
      ADD_u64_u64_408_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : EQ_u16_u1_234_inst 
    ApIntEq_group_15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_0_229;
      iNsTr_1_235 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_234_inst_req_0;
      EQ_u16_u1_234_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_234_inst_req_1;
      EQ_u16_u1_234_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_15_gI: SplitGuardInterface generic map(name => "ApIntEq_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : EQ_u16_u1_386_inst 
    ApIntEq_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rangex_x0_375;
      iNsTr_31_387 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_386_inst_req_0;
      EQ_u16_u1_386_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_386_inst_req_1;
      EQ_u16_u1_386_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_16_gI: SplitGuardInterface generic map(name => "ApIntEq_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : EQ_u16_u1_525_inst 
    ApIntEq_group_17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_44_450 & iNsTr_42_427;
      iNsTr_53_526 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_525_inst_req_0;
      EQ_u16_u1_525_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_525_inst_req_1;
      EQ_u16_u1_525_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_17_gI: SplitGuardInterface generic map(name => "ApIntEq_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : EQ_u16_u1_619_inst 
    ApIntEq_group_18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_55_615 & rangex_x0_375;
      exitcond1_620 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_619_inst_req_0;
      EQ_u16_u1_619_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_619_inst_req_1;
      EQ_u16_u1_619_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_18_gI: SplitGuardInterface generic map(name => "ApIntEq_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : EQ_u16_u1_678_inst 
    ApIntEq_group_19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_674 & rangex_x0_375;
      exitcond_679 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_678_inst_req_0;
      EQ_u16_u1_678_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_678_inst_req_1;
      EQ_u16_u1_678_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_19_gI: SplitGuardInterface generic map(name => "ApIntEq_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : EQ_u32_u1_289_inst 
    ApIntEq_group_20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_9_272 & iNsTr_12_285;
      iNsTr_13_290 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_289_inst_req_0;
      EQ_u32_u1_289_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_289_inst_req_1;
      EQ_u32_u1_289_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_20_gI: SplitGuardInterface generic map(name => "ApIntEq_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : EQ_u8_u1_553_inst 
    ApIntEq_group_21: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= flagx_x12_464;
      iNsTr_59_554 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_553_inst_req_0;
      EQ_u8_u1_553_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_553_inst_req_1;
      EQ_u8_u1_553_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_21_gI: SplitGuardInterface generic map(name => "ApIntEq_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : EQ_u8_u1_641_inst 
    ApIntEq_group_22: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= exorx_x1x_xlcssa_628;
      iNsTr_61_642 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_641_inst_req_0;
      EQ_u8_u1_641_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_641_inst_req_1;
      EQ_u8_u1_641_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_22_gI: SplitGuardInterface generic map(name => "ApIntEq_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : MUL_f32_f32_654_inst 
    ApFloatMul_group_23: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= valx_x1x_xlcssa_632 & signx_x0_650;
      iNsTr_62_655 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= MUL_f32_f32_654_inst_req_0;
      MUL_f32_f32_654_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= MUL_f32_f32_654_inst_req_1;
      MUL_f32_f32_654_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      ApFloatMul_group_23_gI: SplitGuardInterface generic map(name => "ApFloatMul_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatMul_group_23",
          operator_id => "ApFloatMul",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 1,
          use_input_buffering => true,
          full_rate => false,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : SLT_f32_u1_565_inst 
    ApFloatUlt_group_24: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= temp1x_x0_515 & valx_x23_457;
      iNsTr_68_566 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f32_u1_565_inst_req_0;
      SLT_f32_u1_565_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f32_u1_565_inst_req_1;
      SLT_f32_u1_565_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUlt_group_24_gI: SplitGuardInterface generic map(name => "ApFloatUlt_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_24",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : SLT_f64_u1_498_inst 
    ApFloatUlt_group_25: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_48_493;
      iNsTr_49_499 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_498_inst_req_0;
      SLT_f64_u1_498_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_498_inst_req_1;
      SLT_f64_u1_498_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUlt_group_25_gI: SplitGuardInterface generic map(name => "ApFloatUlt_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_25",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : SLT_f64_u1_538_inst 
    ApFloatUlt_group_26: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_48_493;
      iNsTr_57_539 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_538_inst_req_0;
      SLT_f64_u1_538_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_538_inst_req_1;
      SLT_f64_u1_538_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUlt_group_26_gI: SplitGuardInterface generic map(name => "ApFloatUlt_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_26",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : SUB_f32_f32_511_inst 
    ApFloatSub_group_27: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_509_wire_constant & iNsTr_47_489;
      iNsTr_51_512 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_f32_f32_511_inst_req_0;
      SUB_f32_f32_511_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_f32_f32_511_inst_req_1;
      SUB_f32_f32_511_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      ApFloatSub_group_27_gI: SplitGuardInterface generic map(name => "ApFloatSub_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatSub_group_27",
          operator_id => "ApFloatSub",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 1,
          use_input_buffering => true,
          full_rate => false,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : SUB_u16_u16_349_inst 
    ApIntSub_group_28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_28_345 & iNsTr_27_341;
      iNsTr_29_350 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_349_inst_req_0;
      SUB_u16_u16_349_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_349_inst_req_1;
      SUB_u16_u16_349_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_28_gI: SplitGuardInterface generic map(name => "ApIntSub_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : SUB_u16_u16_371_inst 
    ApIntSub_group_29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xneg1_367 & iNsTr_20_361;
      iNsTr_21_372 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_371_inst_req_0;
      SUB_u16_u16_371_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_371_inst_req_1;
      SUB_u16_u16_371_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_29_gI: SplitGuardInterface generic map(name => "ApIntSub_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : ULT_u16_u1_692_inst 
    ApIntUlt_group_30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp17_258 & iNsTr_10_275;
      iNsTr_33_693 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u16_u1_692_inst_req_0;
      ULT_u16_u1_692_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u16_u1_692_inst_req_1;
      ULT_u16_u1_692_inst_ack_1 <= ackR_unguarded(0);
      ApIntUlt_group_30_gI: SplitGuardInterface generic map(name => "ApIntUlt_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : XOR_u8_u8_547_inst 
    ApIntXor_group_31: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_58_543 & exorx_x25_442;
      exorx_x0_548 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u8_u8_547_inst_req_0;
      XOR_u8_u8_547_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u8_u8_547_inst_req_1;
      XOR_u8_u8_547_inst_ack_1 <= ackR_unguarded(0);
      ApIntXor_group_31_gI: SplitGuardInterface generic map(name => "ApIntXor_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : type_cast_492_inst 
    ApFloatResize_group_32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_47_489;
      iNsTr_48_493 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_492_inst_req_0;
      type_cast_492_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_492_inst_req_1;
      type_cast_492_inst_ack_1 <= ackR_unguarded(0);
      ApFloatResize_group_32_gI: SplitGuardInterface generic map(name => "ApFloatResize_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApFloatResize_group_32",
          operator_id => "ApFloatResize",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 1,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : LOAD_ncol_ind_266_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_ncol_ind_266_load_0_req_0;
      LOAD_ncol_ind_266_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ncol_ind_266_load_0_req_1;
      LOAD_ncol_ind_266_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncol_ind_266_word_address_0;
      LOAD_ncol_ind_266_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(15 downto 0),
          mtag => memory_space_10_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_nrows_274_load_0 LOAD_nrows_228_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= LOAD_nrows_274_load_0_req_0;
      reqL_unguarded(0) <= LOAD_nrows_228_load_0_req_0;
      LOAD_nrows_274_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_nrows_228_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_nrows_274_load_0_req_1;
      reqR_unguarded(0) <= LOAD_nrows_228_load_0_req_1;
      LOAD_nrows_274_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_nrows_228_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_nrows_274_word_address_0 & LOAD_nrows_228_word_address_0;
      LOAD_nrows_274_data_0 <= data_out(31 downto 16);
      LOAD_nrows_228_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_12_lr_req(0),
          mack => memory_space_12_lr_ack(0),
          maddr => memory_space_12_lr_addr(0 downto 0),
          mtag => memory_space_12_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_12_lc_req(0),
          mack => memory_space_12_lc_ack(0),
          mdata => memory_space_12_lc_data(15 downto 0),
          mtag => memory_space_12_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_340_load_0 ptr_deref_417_load_0 ptr_deref_360_load_0 ptr_deref_344_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_340_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_417_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_360_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_344_load_0_req_0;
      ptr_deref_340_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_417_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_360_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_344_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_340_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_417_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_360_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_344_load_0_req_1;
      ptr_deref_340_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_417_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_360_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_344_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_340_word_address_0 & ptr_deref_417_word_address_0 & ptr_deref_360_word_address_0 & ptr_deref_344_word_address_0;
      ptr_deref_340_data_0 <= data_out(63 downto 48);
      ptr_deref_417_data_0 <= data_out(47 downto 32);
      ptr_deref_360_data_0 <= data_out(31 downto 16);
      ptr_deref_344_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 10,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(9 downto 0),
          mtag => memory_space_8_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_488_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_488_load_0_req_0;
      ptr_deref_488_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_488_load_0_req_1;
      ptr_deref_488_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_488_word_address_0;
      ptr_deref_488_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 10,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(9 downto 0),
          mtag => memory_space_9_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(31 downto 0),
          mtag => memory_space_9_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_666_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_666_store_0_req_0;
      ptr_deref_666_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_666_store_0_req_1;
      ptr_deref_666_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_666_word_address_0;
      data_in <= ptr_deref_666_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(9 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end checkNodeComputeEngine_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity initInputs is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_11_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_11_sr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_10_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_12_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_12_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_12_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_12_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_12_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_12_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_13_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_13_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_13_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_13_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_13_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_13_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_sc_tag :  in  std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    matrix_in_pipe_read_req : out  std_logic_vector(1 downto 0);
    matrix_in_pipe_read_ack : in   std_logic_vector(1 downto 0);
    matrix_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
    rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initInputs;
architecture initInputs_arch of initInputs is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal initInputs_CP_3524_start: Boolean;
  signal initInputs_CP_3524_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal STORE_nrows_793_store_0_ack_0 : boolean;
  signal ADD_u64_u64_768_inst_req_0 : boolean;
  signal ptr_deref_761_store_0_ack_0 : boolean;
  signal ptr_deref_761_store_0_req_0 : boolean;
  signal EQ_u64_u1_774_inst_req_0 : boolean;
  signal ADD_u64_u64_768_inst_ack_1 : boolean;
  signal ADD_u64_u64_768_inst_req_1 : boolean;
  signal STORE_nrows_793_store_0_req_0 : boolean;
  signal ptr_deref_761_store_0_ack_1 : boolean;
  signal ptr_deref_791_load_0_ack_1 : boolean;
  signal EQ_u64_u1_774_inst_ack_0 : boolean;
  signal ADD_u64_u64_768_inst_ack_0 : boolean;
  signal ptr_deref_761_store_0_req_1 : boolean;
  signal STORE_nrows_793_store_0_req_1 : boolean;
  signal STORE_nrows_793_store_0_ack_1 : boolean;
  signal ptr_deref_791_load_0_req_1 : boolean;
  signal if_stmt_776_branch_ack_0 : boolean;
  signal STORE_ncols_806_store_0_req_0 : boolean;
  signal STORE_ncols_806_store_0_ack_0 : boolean;
  signal ptr_deref_804_load_0_req_1 : boolean;
  signal ptr_deref_804_load_0_ack_1 : boolean;
  signal ptr_deref_804_load_0_req_0 : boolean;
  signal ptr_deref_804_load_0_ack_0 : boolean;
  signal STORE_ncols_806_store_0_req_1 : boolean;
  signal STORE_ncols_806_store_0_ack_1 : boolean;
  signal if_stmt_776_branch_ack_1 : boolean;
  signal ptr_deref_791_load_0_ack_0 : boolean;
  signal ptr_deref_791_load_0_req_0 : boolean;
  signal if_stmt_776_branch_req_0 : boolean;
  signal EQ_u64_u1_774_inst_ack_1 : boolean;
  signal EQ_u64_u1_774_inst_req_1 : boolean;
  signal RPIPE_maxNitr_in_731_inst_req_0 : boolean;
  signal RPIPE_maxNitr_in_731_inst_ack_0 : boolean;
  signal RPIPE_maxNitr_in_731_inst_req_1 : boolean;
  signal RPIPE_maxNitr_in_731_inst_ack_1 : boolean;
  signal STORE_maxNitr_733_store_0_req_0 : boolean;
  signal STORE_maxNitr_733_store_0_ack_0 : boolean;
  signal STORE_maxNitr_733_store_0_req_1 : boolean;
  signal STORE_maxNitr_733_store_0_ack_1 : boolean;
  signal RPIPE_ebbyNo_in_737_inst_req_0 : boolean;
  signal RPIPE_ebbyNo_in_737_inst_ack_0 : boolean;
  signal RPIPE_ebbyNo_in_737_inst_req_1 : boolean;
  signal RPIPE_ebbyNo_in_737_inst_ack_1 : boolean;
  signal STORE_ebbyNo_739_store_0_req_0 : boolean;
  signal STORE_ebbyNo_739_store_0_ack_0 : boolean;
  signal STORE_ebbyNo_739_store_0_req_1 : boolean;
  signal STORE_ebbyNo_739_store_0_ack_1 : boolean;
  signal addr_of_755_final_reg_req_0 : boolean;
  signal addr_of_755_final_reg_ack_0 : boolean;
  signal addr_of_755_final_reg_req_1 : boolean;
  signal addr_of_755_final_reg_ack_1 : boolean;
  signal RPIPE_matrix_in_758_inst_req_0 : boolean;
  signal RPIPE_matrix_in_758_inst_ack_0 : boolean;
  signal RPIPE_matrix_in_758_inst_req_1 : boolean;
  signal RPIPE_matrix_in_758_inst_ack_1 : boolean;
  signal ptr_deref_817_load_0_req_0 : boolean;
  signal ptr_deref_817_load_0_ack_0 : boolean;
  signal ptr_deref_817_load_0_req_1 : boolean;
  signal ptr_deref_817_load_0_ack_1 : boolean;
  signal STORE_ncol_ind_819_store_0_req_0 : boolean;
  signal STORE_ncol_ind_819_store_0_ack_0 : boolean;
  signal STORE_ncol_ind_819_store_0_req_1 : boolean;
  signal STORE_ncol_ind_819_store_0_ack_1 : boolean;
  signal SUB_u16_u16_826_inst_req_0 : boolean;
  signal SUB_u16_u16_826_inst_ack_0 : boolean;
  signal SUB_u16_u16_826_inst_req_1 : boolean;
  signal SUB_u16_u16_826_inst_ack_1 : boolean;
  signal EQ_u16_u1_831_inst_req_0 : boolean;
  signal EQ_u16_u1_831_inst_ack_0 : boolean;
  signal EQ_u16_u1_831_inst_req_1 : boolean;
  signal EQ_u16_u1_831_inst_ack_1 : boolean;
  signal if_stmt_833_branch_req_0 : boolean;
  signal if_stmt_833_branch_ack_1 : boolean;
  signal if_stmt_833_branch_ack_0 : boolean;
  signal ADD_u16_u16_843_inst_req_0 : boolean;
  signal ADD_u16_u16_843_inst_ack_0 : boolean;
  signal ADD_u16_u16_843_inst_req_1 : boolean;
  signal ADD_u16_u16_843_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal do_while_stmt_857_branch_req_0 : boolean;
  signal phi_stmt_859_req_0 : boolean;
  signal phi_stmt_859_req_1 : boolean;
  signal phi_stmt_859_ack_0 : boolean;
  signal type_cast_862_inst_req_0 : boolean;
  signal type_cast_862_inst_ack_0 : boolean;
  signal type_cast_862_inst_req_1 : boolean;
  signal type_cast_862_inst_ack_1 : boolean;
  signal indvar_at_entry_851_863_buf_req_0 : boolean;
  signal indvar_at_entry_851_863_buf_ack_0 : boolean;
  signal indvar_at_entry_851_863_buf_req_1 : boolean;
  signal indvar_at_entry_851_863_buf_ack_1 : boolean;
  signal ADD_u64_u64_869_inst_req_0 : boolean;
  signal ADD_u64_u64_869_inst_ack_0 : boolean;
  signal ADD_u64_u64_869_inst_req_1 : boolean;
  signal ADD_u64_u64_869_inst_ack_1 : boolean;
  signal addr_of_874_final_reg_req_0 : boolean;
  signal addr_of_874_final_reg_ack_0 : boolean;
  signal addr_of_874_final_reg_req_1 : boolean;
  signal addr_of_874_final_reg_ack_1 : boolean;
  signal RPIPE_matrix_in_877_inst_req_0 : boolean;
  signal RPIPE_matrix_in_877_inst_ack_0 : boolean;
  signal RPIPE_matrix_in_877_inst_req_1 : boolean;
  signal RPIPE_matrix_in_877_inst_ack_1 : boolean;
  signal ptr_deref_880_store_0_req_0 : boolean;
  signal ptr_deref_880_store_0_ack_0 : boolean;
  signal ptr_deref_880_store_0_req_1 : boolean;
  signal ptr_deref_880_store_0_ack_1 : boolean;
  signal ADD_u64_u64_887_inst_req_0 : boolean;
  signal ADD_u64_u64_887_inst_ack_0 : boolean;
  signal ADD_u64_u64_887_inst_req_1 : boolean;
  signal ADD_u64_u64_887_inst_ack_1 : boolean;
  signal EQ_u64_u1_892_inst_req_0 : boolean;
  signal EQ_u64_u1_892_inst_ack_0 : boolean;
  signal EQ_u64_u1_892_inst_req_1 : boolean;
  signal EQ_u64_u1_892_inst_ack_1 : boolean;
  signal W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_0 : boolean;
  signal W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_0 : boolean;
  signal W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_1 : boolean;
  signal W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_1 : boolean;
  signal do_while_stmt_857_branch_ack_0 : boolean;
  signal do_while_stmt_857_branch_ack_1 : boolean;
  signal if_stmt_900_branch_req_0 : boolean;
  signal if_stmt_900_branch_ack_1 : boolean;
  signal if_stmt_900_branch_ack_0 : boolean;
  signal RPIPE_rate_in_908_inst_req_0 : boolean;
  signal RPIPE_rate_in_908_inst_ack_0 : boolean;
  signal RPIPE_rate_in_908_inst_req_1 : boolean;
  signal RPIPE_rate_in_908_inst_ack_1 : boolean;
  signal STORE_rate_910_store_0_req_0 : boolean;
  signal STORE_rate_910_store_0_ack_0 : boolean;
  signal STORE_rate_910_store_0_req_1 : boolean;
  signal STORE_rate_910_store_0_ack_1 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal phi_stmt_744_req_1 : boolean;
  signal phi_stmt_744_req_0 : boolean;
  signal phi_stmt_744_ack_0 : boolean;
  signal phi_stmt_851_req_0 : boolean;
  signal phi_stmt_851_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initInputs_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initInputs_CP_3524_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initInputs_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initInputs_CP_3524_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initInputs_CP_3524_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initInputs_CP_3524_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initInputs_CP_3524: Block -- control-path 
    signal initInputs_CP_3524_elements: BooleanArray(208 downto 0);
    -- 
  begin -- 
    initInputs_CP_3524_elements(0) <= initInputs_CP_3524_start;
    initInputs_CP_3524_symbol <= initInputs_CP_3524_elements(207);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_729/$entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	22 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_729/branch_block_stmt_729__entry__
      -- CP-element group 1: 	 branch_block_stmt_729/assign_stmt_732__entry__
      -- 
    initInputs_CP_3524_elements(1) <= initInputs_CP_3524_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	24 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	25 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_729/assign_stmt_732__exit__
      -- CP-element group 2: 	 branch_block_stmt_729/assign_stmt_735__entry__
      -- 
    initInputs_CP_3524_elements(2) <= initInputs_CP_3524_elements(24);
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	27 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_729/assign_stmt_735__exit__
      -- CP-element group 3: 	 branch_block_stmt_729/assign_stmt_738__entry__
      -- 
    initInputs_CP_3524_elements(3) <= initInputs_CP_3524_elements(27);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	30 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	31 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_729/assign_stmt_738__exit__
      -- CP-element group 4: 	 branch_block_stmt_729/assign_stmt_741__entry__
      -- 
    initInputs_CP_3524_elements(4) <= initInputs_CP_3524_elements(30);
    -- CP-element group 5:  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	33 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	178 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_729/assign_stmt_741__exit__
      -- CP-element group 5: 	 branch_block_stmt_729/bbx_xnph3_bb_1
      -- 
    initInputs_CP_3524_elements(5) <= initInputs_CP_3524_elements(33);
    -- CP-element group 6:  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	183 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	34 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_729/merge_stmt_743__exit__
      -- CP-element group 6: 	 branch_block_stmt_729/assign_stmt_756__entry__
      -- 
    initInputs_CP_3524_elements(6) <= initInputs_CP_3524_elements(183);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	37 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	38 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_729/assign_stmt_756__exit__
      -- CP-element group 7: 	 branch_block_stmt_729/assign_stmt_759__entry__
      -- 
    initInputs_CP_3524_elements(7) <= initInputs_CP_3524_elements(37);
    -- CP-element group 8:  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	40 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	41 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_729/assign_stmt_759__exit__
      -- CP-element group 8: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775__entry__
      -- 
    initInputs_CP_3524_elements(8) <= initInputs_CP_3524_elements(40);
    -- CP-element group 9:  branch  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	48 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	49 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775__exit__
      -- CP-element group 9: 	 branch_block_stmt_729/if_stmt_776__entry__
      -- 
    initInputs_CP_3524_elements(9) <= initInputs_CP_3524_elements(48);
    -- CP-element group 10:  merge  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	186 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	58 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_729/merge_stmt_782__exit__
      -- CP-element group 10: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832__entry__
      -- 
    initInputs_CP_3524_elements(10) <= initInputs_CP_3524_elements(186);
    -- CP-element group 11:  branch  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	79 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	80 
    -- CP-element group 11: 	81 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832__exit__
      -- CP-element group 11: 	 branch_block_stmt_729/if_stmt_833__entry__
      -- 
    initInputs_CP_3524_elements(11) <= initInputs_CP_3524_elements(79);
    -- CP-element group 12:  merge  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	189 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	89 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_729/merge_stmt_839__exit__
      -- CP-element group 12: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848__entry__
      -- 
    initInputs_CP_3524_elements(12) <= initInputs_CP_3524_elements(189);
    -- CP-element group 13:  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	93 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	190 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848__exit__
      -- CP-element group 13: 	 branch_block_stmt_729/bbx_xnph_bb_4
      -- 
    initInputs_CP_3524_elements(13) <= initInputs_CP_3524_elements(93);
    -- CP-element group 14:  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	195 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	94 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_729/merge_stmt_850__exit__
      -- CP-element group 14: 	 branch_block_stmt_729/do_while_stmt_857__entry__
      -- 
    initInputs_CP_3524_elements(14) <= initInputs_CP_3524_elements(195);
    -- CP-element group 15:  branch  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	159 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	160 
    -- CP-element group 15: 	161 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_729/do_while_stmt_857__exit__
      -- CP-element group 15: 	 branch_block_stmt_729/if_stmt_900__entry__
      -- 
    initInputs_CP_3524_elements(15) <= initInputs_CP_3524_elements(159);
    -- CP-element group 16:  merge  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	166 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	196 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_729/if_stmt_900__exit__
      -- CP-element group 16: 	 branch_block_stmt_729/merge_stmt_904__entry__
      -- 
    initInputs_CP_3524_elements(16) <= initInputs_CP_3524_elements(166);
    -- CP-element group 17:  merge  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	199 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	201 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_729/merge_stmt_904__exit__
      -- CP-element group 17: 	 branch_block_stmt_729/xx_x_crit_edgex_xloopexit_xx_x_crit_edge
      -- 
    initInputs_CP_3524_elements(17) <= initInputs_CP_3524_elements(199);
    -- CP-element group 18:  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	203 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	168 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_729/merge_stmt_906__exit__
      -- CP-element group 18: 	 branch_block_stmt_729/assign_stmt_909__entry__
      -- 
    initInputs_CP_3524_elements(18) <= initInputs_CP_3524_elements(203);
    -- CP-element group 19:  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	170 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	171 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_729/assign_stmt_909__exit__
      -- CP-element group 19: 	 branch_block_stmt_729/assign_stmt_912__entry__
      -- 
    initInputs_CP_3524_elements(19) <= initInputs_CP_3524_elements(170);
    -- CP-element group 20:  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	173 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	204 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_729/assign_stmt_912__exit__
      -- CP-element group 20: 	 branch_block_stmt_729/return__
      -- 
    initInputs_CP_3524_elements(20) <= initInputs_CP_3524_elements(173);
    -- CP-element group 21:  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	206 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	207 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_729/branch_block_stmt_729__exit__
      -- CP-element group 21: 	 branch_block_stmt_729/merge_stmt_914__exit__
      -- 
    initInputs_CP_3524_elements(21) <= initInputs_CP_3524_elements(206);
    -- CP-element group 22:  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_729/assign_stmt_732/$entry
      -- CP-element group 22: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Sample/rr
      -- 
    rr_3586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(22), ack => RPIPE_maxNitr_in_731_inst_req_0); -- 
    initInputs_CP_3524_elements(22) <= initInputs_CP_3524_elements(1);
    -- CP-element group 23:  transition  input  output  no-bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_update_start_
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Update/cr
      -- 
    ra_3587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxNitr_in_731_inst_ack_0, ack => initInputs_CP_3524_elements(23)); -- 
    cr_3591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(23), ack => RPIPE_maxNitr_in_731_inst_req_1); -- 
    -- CP-element group 24:  transition  input  no-bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	2 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_729/assign_stmt_732/$exit
      -- CP-element group 24: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_729/assign_stmt_732/RPIPE_maxNitr_in_731_Update/ca
      -- 
    ca_3592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxNitr_in_731_inst_ack_1, ack => initInputs_CP_3524_elements(24)); -- 
    -- CP-element group 25:  fork  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (17) 
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_update_start_
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_word_address_calculated
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_root_address_calculated
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/STORE_maxNitr_733_Split/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/STORE_maxNitr_733_Split/$exit
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/STORE_maxNitr_733_Split/split_req
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/STORE_maxNitr_733_Split/split_ack
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/word_0/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/word_0/rr
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/word_0/$entry
      -- CP-element group 25: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/word_0/cr
      -- 
    cr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(25), ack => STORE_maxNitr_733_store_0_req_1); -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(25), ack => STORE_maxNitr_733_store_0_req_0); -- 
    initInputs_CP_3524_elements(25) <= initInputs_CP_3524_elements(2);
    -- CP-element group 26:  transition  input  no-bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/$exit
      -- CP-element group 26: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Sample/word_access_start/word_0/ra
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_maxNitr_733_store_0_ack_0, ack => initInputs_CP_3524_elements(26)); -- 
    -- CP-element group 27:  transition  input  no-bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	3 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/$exit
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/$exit
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_729/assign_stmt_735/STORE_maxNitr_733_Update/word_access_complete/word_0/ca
      -- 
    ca_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_maxNitr_733_store_0_ack_1, ack => initInputs_CP_3524_elements(27)); -- 
    -- CP-element group 28:  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_729/assign_stmt_738/$entry
      -- CP-element group 28: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Sample/rr
      -- 
    rr_3639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(28), ack => RPIPE_ebbyNo_in_737_inst_req_0); -- 
    initInputs_CP_3524_elements(28) <= initInputs_CP_3524_elements(3);
    -- CP-element group 29:  transition  input  output  no-bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_update_start_
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Update/cr
      -- 
    ra_3640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ebbyNo_in_737_inst_ack_0, ack => initInputs_CP_3524_elements(29)); -- 
    cr_3644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(29), ack => RPIPE_ebbyNo_in_737_inst_req_1); -- 
    -- CP-element group 30:  transition  input  no-bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	4 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_729/assign_stmt_738/$exit
      -- CP-element group 30: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_729/assign_stmt_738/RPIPE_ebbyNo_in_737_Update/ca
      -- 
    ca_3645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ebbyNo_in_737_inst_ack_1, ack => initInputs_CP_3524_elements(30)); -- 
    -- CP-element group 31:  fork  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	4 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (17) 
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_update_start_
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/STORE_ebbyNo_739_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/STORE_ebbyNo_739_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/STORE_ebbyNo_739_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/STORE_ebbyNo_739_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/word_0/cr
      -- 
    cr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(31), ack => STORE_ebbyNo_739_store_0_req_1); -- 
    rr_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(31), ack => STORE_ebbyNo_739_store_0_req_0); -- 
    initInputs_CP_3524_elements(31) <= initInputs_CP_3524_elements(4);
    -- CP-element group 32:  transition  input  no-bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Sample/word_access_start/word_0/ra
      -- 
    ra_3670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ebbyNo_739_store_0_ack_0, ack => initInputs_CP_3524_elements(32)); -- 
    -- CP-element group 33:  transition  input  no-bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	5 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/$exit
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_729/assign_stmt_741/STORE_ebbyNo_739_Update/word_access_complete/word_0/ca
      -- 
    ca_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ebbyNo_739_store_0_ack_1, ack => initInputs_CP_3524_elements(33)); -- 
    -- CP-element group 34:  fork  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	6 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_update_start_
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_root_address_calculated
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_offset_calculated
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_resized_0
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_scaled_0
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_computed_0
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_resize_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_resize_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_resize_0/index_resize_req
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_resize_0/index_resize_ack
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_scale_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_scale_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_scale_0/scale_rename_req
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_index_scale_0/scale_rename_ack
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_final_index_sum_regn/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_final_index_sum_regn/$exit
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_final_index_sum_regn/req
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_final_index_sum_regn/ack
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_base_plus_offset/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_base_plus_offset/$exit
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_base_plus_offset/sum_rename_req
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/array_obj_ref_754_base_plus_offset/sum_rename_ack
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_request/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_request/req
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_complete/req
      -- 
    req_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(34), ack => addr_of_755_final_reg_req_1); -- 
    req_3717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(34), ack => addr_of_755_final_reg_req_0); -- 
    initInputs_CP_3524_elements(34) <= initInputs_CP_3524_elements(6);
    -- CP-element group 35:  transition  input  no-bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_request/$exit
      -- CP-element group 35: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_request/ack
      -- 
    ack_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_755_final_reg_ack_0, ack => initInputs_CP_3524_elements(35)); -- 
    -- CP-element group 36:  transition  input  no-bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_729/assign_stmt_756/addr_of_755_complete/ack
      -- 
    ack_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_755_final_reg_ack_1, ack => initInputs_CP_3524_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	7 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_729/assign_stmt_756/$exit
      -- 
    initInputs_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(35) & initInputs_CP_3524_elements(36);
      gj_initInputs_cp_element_group_37 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_729/assign_stmt_759/$entry
      -- CP-element group 38: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Sample/rr
      -- 
    rr_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(38), ack => RPIPE_matrix_in_758_inst_req_0); -- 
    initInputs_CP_3524_elements(38) <= initInputs_CP_3524_elements(7);
    -- CP-element group 39:  transition  input  output  no-bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_update_start_
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Update/cr
      -- 
    ra_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_758_inst_ack_0, ack => initInputs_CP_3524_elements(39)); -- 
    cr_3739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(39), ack => RPIPE_matrix_in_758_inst_req_1); -- 
    -- CP-element group 40:  transition  input  no-bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	8 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_729/assign_stmt_759/$exit
      -- CP-element group 40: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_729/assign_stmt_759/RPIPE_matrix_in_758_Update/ca
      -- 
    ca_3740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_758_inst_ack_1, ack => initInputs_CP_3524_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	8 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	44 
    -- CP-element group 41: 	45 
    -- CP-element group 41: 	47 
    -- CP-element group 41:  members (40) 
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/ptr_deref_761_Split/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/ptr_deref_761_Split/split_ack
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_update_start_
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/ptr_deref_761_Split/split_req
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/ptr_deref_761_Split/$exit
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_update_start_
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/$entry
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_update_start_
      -- CP-element group 41: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_base_address_calculated
      -- 
    cr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(41), ack => ptr_deref_761_store_0_req_1); -- 
    rr_3781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(41), ack => ptr_deref_761_store_0_req_0); -- 
    rr_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(41), ack => ADD_u64_u64_768_inst_req_0); -- 
    cr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(41), ack => ADD_u64_u64_768_inst_req_1); -- 
    cr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(41), ack => EQ_u64_u1_774_inst_req_1); -- 
    initInputs_CP_3524_elements(41) <= initInputs_CP_3524_elements(8);
    -- CP-element group 42:  transition  input  no-bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/word_0/ra
      -- CP-element group 42: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_sample_completed_
      -- 
    ra_3782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_761_store_0_ack_0, ack => initInputs_CP_3524_elements(42)); -- 
    -- CP-element group 43:  transition  input  no-bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ptr_deref_761_update_completed_
      -- 
    ca_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_761_store_0_ack_1, ack => initInputs_CP_3524_elements(43)); -- 
    -- CP-element group 44:  transition  input  no-bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	41 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_sample_completed_
      -- 
    ra_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_768_inst_ack_0, ack => initInputs_CP_3524_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  no-bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	41 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/ADD_u64_u64_768_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Sample/$entry
      -- 
    ca_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_768_inst_ack_1, ack => initInputs_CP_3524_elements(45)); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(45), ack => EQ_u64_u1_774_inst_req_0); -- 
    -- CP-element group 46:  transition  input  no-bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Sample/ra
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_774_inst_ack_0, ack => initInputs_CP_3524_elements(46)); -- 
    -- CP-element group 47:  transition  input  no-bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	41 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/EQ_u64_u1_774_Update/$exit
      -- 
    ca_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_774_inst_ack_1, ack => initInputs_CP_3524_elements(47)); -- 
    -- CP-element group 48:  join  transition  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	9 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_729/assign_stmt_763_to_assign_stmt_775/$exit
      -- 
    initInputs_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(43) & initInputs_CP_3524_elements(47);
      gj_initInputs_cp_element_group_48 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	9 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_729/if_stmt_776_dead_link/$entry
      -- 
    initInputs_CP_3524_elements(49) <= initInputs_CP_3524_elements(9);
    -- CP-element group 50:  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	9 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_729/if_stmt_776_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_729/if_stmt_776_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_729/if_stmt_776_eval_test/$entry
      -- 
    branch_req_3829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(50), ack => if_stmt_776_branch_req_0); -- 
    initInputs_CP_3524_elements(50) <= initInputs_CP_3524_elements(9);
    -- CP-element group 51:  branch  place  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_729/R_exitcond_777_place
      -- 
    initInputs_CP_3524_elements(51) <= initInputs_CP_3524_elements(50);
    -- CP-element group 52:  transition  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_729/if_stmt_776_if_link/$entry
      -- 
    initInputs_CP_3524_elements(52) <= initInputs_CP_3524_elements(51);
    -- CP-element group 53:  transition  input  no-bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_729/if_stmt_776_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_729/if_stmt_776_if_link/$exit
      -- 
    if_choice_transition_3834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_776_branch_ack_1, ack => initInputs_CP_3524_elements(53)); -- 
    -- CP-element group 54:  transition  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_729/if_stmt_776_else_link/$entry
      -- 
    initInputs_CP_3524_elements(54) <= initInputs_CP_3524_elements(51);
    -- CP-element group 55:  transition  input  no-bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_729/if_stmt_776_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_729/if_stmt_776_else_link/$exit
      -- 
    else_choice_transition_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_776_branch_ack_0, ack => initInputs_CP_3524_elements(55)); -- 
    -- CP-element group 56:  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	184 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_729/bb_1_xx_x_crit_edge4
      -- 
    initInputs_CP_3524_elements(56) <= initInputs_CP_3524_elements(53);
    -- CP-element group 57:  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	174 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_729/bb_1_bb_1
      -- 
    initInputs_CP_3524_elements(57) <= initInputs_CP_3524_elements(55);
    -- CP-element group 58:  join  fork  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	10 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	61 
    -- CP-element group 58: 	63 
    -- CP-element group 58: 	64 
    -- CP-element group 58: 	65 
    -- CP-element group 58: 	66 
    -- CP-element group 58: 	68 
    -- CP-element group 58: 	69 
    -- CP-element group 58: 	70 
    -- CP-element group 58: 	71 
    -- CP-element group 58: 	73 
    -- CP-element group 58: 	75 
    -- CP-element group 58: 	78 
    -- CP-element group 58:  members (106) 
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/word_0/rr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/word_0/rr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/word_0/rr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_update_start_
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Update/cr
      -- 
    cr_3887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_791_load_0_req_1); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_791_load_0_req_0); -- 
    cr_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => STORE_nrows_793_store_0_req_1); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_804_load_0_req_1); -- 
    rr_3959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_804_load_0_req_0); -- 
    cr_4008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => STORE_ncols_806_store_0_req_1); -- 
    cr_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_817_load_0_req_1); -- 
    rr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => ptr_deref_817_load_0_req_0); -- 
    cr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => STORE_ncol_ind_819_store_0_req_1); -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => SUB_u16_u16_826_inst_req_1); -- 
    cr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(58), ack => EQ_u16_u1_831_inst_req_1); -- 
    initInputs_CP_3524_elements(58) <= initInputs_CP_3524_elements(10);
    -- CP-element group 59:  transition  input  no-bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/word_0/ra
      -- CP-element group 59: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Sample/word_access_start/word_0/$exit
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_791_load_0_ack_0, ack => initInputs_CP_3524_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  no-bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	76 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/ptr_deref_791_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/ptr_deref_791_Merge/merge_ack
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/ptr_deref_791_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/ptr_deref_791_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_791_Update/$exit
      -- 
    ca_3888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_791_load_0_ack_1, ack => initInputs_CP_3524_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  no-bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/STORE_nrows_793_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/word_0/rr
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/STORE_nrows_793_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/STORE_nrows_793_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/STORE_nrows_793_Split/$entry
      -- 
    rr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(61), ack => STORE_nrows_793_store_0_req_0); -- 
    initInputs_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(58) & initInputs_CP_3524_elements(60);
      gj_initInputs_cp_element_group_61 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  no-bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/word_0/ra
      -- CP-element group 62: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Sample/$exit
      -- 
    ra_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_nrows_793_store_0_ack_0, ack => initInputs_CP_3524_elements(62)); -- 
    -- CP-element group 63:  transition  input  no-bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	58 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	79 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/word_0/ca
      -- CP-element group 63: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_nrows_793_Update/word_access_complete/word_0/$exit
      -- 
    ca_3926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_nrows_793_store_0_ack_1, ack => initInputs_CP_3524_elements(63)); -- 
    -- CP-element group 64:  transition  input  no-bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Sample/word_access_start/word_0/ra
      -- 
    ra_3960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_804_load_0_ack_0, ack => initInputs_CP_3524_elements(64)); -- 
    -- CP-element group 65:  transition  input  no-bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	58 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (9) 
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/ptr_deref_804_Merge/$entry
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/ptr_deref_804_Merge/$exit
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/ptr_deref_804_Merge/merge_req
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_804_Update/ptr_deref_804_Merge/merge_ack
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_804_load_0_ack_1, ack => initInputs_CP_3524_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  no-bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	58 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/$entry
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/word_0/$entry
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/STORE_ncols_806_Split/$entry
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/STORE_ncols_806_Split/$exit
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/STORE_ncols_806_Split/split_req
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/STORE_ncols_806_Split/split_ack
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/word_0/rr
      -- 
    rr_3997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(66), ack => STORE_ncols_806_store_0_req_0); -- 
    initInputs_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(58) & initInputs_CP_3524_elements(65);
      gj_initInputs_cp_element_group_66 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  no-bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/$exit
      -- CP-element group 67: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/word_0/$exit
      -- CP-element group 67: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Sample/word_access_start/word_0/ra
      -- 
    ra_3998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncols_806_store_0_ack_0, ack => initInputs_CP_3524_elements(67)); -- 
    -- CP-element group 68:  transition  input  no-bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	58 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	79 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/$exit
      -- CP-element group 68: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncols_806_Update/word_access_complete/word_0/ca
      -- 
    ca_4009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncols_806_store_0_ack_1, ack => initInputs_CP_3524_elements(68)); -- 
    -- CP-element group 69:  transition  input  no-bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	58 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/$exit
      -- CP-element group 69: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Sample/word_access_start/word_0/ra
      -- 
    ra_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_817_load_0_ack_0, ack => initInputs_CP_3524_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  output  no-bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	58 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (12) 
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/word_access_complete/word_0/ca
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/ptr_deref_817_Merge/$entry
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/ptr_deref_817_Merge/$exit
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/ptr_deref_817_Merge/merge_req
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/ptr_deref_817_Update/ptr_deref_817_Merge/merge_ack
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Sample/rr
      -- 
    ca_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_817_load_0_ack_1, ack => initInputs_CP_3524_elements(70)); -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(70), ack => SUB_u16_u16_826_inst_req_0); -- 
    -- CP-element group 71:  join  transition  output  no-bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	58 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/STORE_ncol_ind_819_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/STORE_ncol_ind_819_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/STORE_ncol_ind_819_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/STORE_ncol_ind_819_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/word_0/rr
      -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(71), ack => STORE_ncol_ind_819_store_0_req_0); -- 
    initInputs_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(58) & initInputs_CP_3524_elements(70);
      gj_initInputs_cp_element_group_71 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  no-bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Sample/word_access_start/word_0/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncol_ind_819_store_0_ack_0, ack => initInputs_CP_3524_elements(72)); -- 
    -- CP-element group 73:  transition  input  no-bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	58 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	79 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/STORE_ncol_ind_819_Update/word_access_complete/word_0/ca
      -- 
    ca_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ncol_ind_819_store_0_ack_1, ack => initInputs_CP_3524_elements(73)); -- 
    -- CP-element group 74:  transition  input  no-bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Sample/ra
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_826_inst_ack_0, ack => initInputs_CP_3524_elements(74)); -- 
    -- CP-element group 75:  transition  input  no-bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	58 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/SUB_u16_u16_826_Update/ca
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_826_inst_ack_1, ack => initInputs_CP_3524_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	60 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Sample/rr
      -- 
    rr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(76), ack => EQ_u16_u1_831_inst_req_0); -- 
    initInputs_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(60) & initInputs_CP_3524_elements(75);
      gj_initInputs_cp_element_group_76 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  no-bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Sample/ra
      -- 
    ra_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_831_inst_ack_0, ack => initInputs_CP_3524_elements(77)); -- 
    -- CP-element group 78:  transition  input  no-bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	58 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/EQ_u16_u1_831_Update/ca
      -- 
    ca_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_831_inst_ack_1, ack => initInputs_CP_3524_elements(78)); -- 
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	63 
    -- CP-element group 79: 	68 
    -- CP-element group 79: 	73 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	11 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_729/assign_stmt_788_to_assign_stmt_832/$exit
      -- 
    initInputs_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "initInputs_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(63) & initInputs_CP_3524_elements(68) & initInputs_CP_3524_elements(73) & initInputs_CP_3524_elements(78);
      gj_initInputs_cp_element_group_79 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	11 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_729/if_stmt_833_dead_link/$entry
      -- 
    initInputs_CP_3524_elements(80) <= initInputs_CP_3524_elements(11);
    -- CP-element group 81:  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	11 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_729/if_stmt_833_eval_test/$entry
      -- CP-element group 81: 	 branch_block_stmt_729/if_stmt_833_eval_test/$exit
      -- CP-element group 81: 	 branch_block_stmt_729/if_stmt_833_eval_test/branch_req
      -- 
    branch_req_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(81), ack => if_stmt_833_branch_req_0); -- 
    initInputs_CP_3524_elements(81) <= initInputs_CP_3524_elements(11);
    -- CP-element group 82:  branch  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_729/R_iNsTr_21_834_place
      -- 
    initInputs_CP_3524_elements(82) <= initInputs_CP_3524_elements(81);
    -- CP-element group 83:  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_729/if_stmt_833_if_link/$entry
      -- 
    initInputs_CP_3524_elements(83) <= initInputs_CP_3524_elements(82);
    -- CP-element group 84:  transition  input  no-bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	87 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_729/if_stmt_833_if_link/$exit
      -- CP-element group 84: 	 branch_block_stmt_729/if_stmt_833_if_link/if_choice_transition
      -- 
    if_choice_transition_4133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_833_branch_ack_1, ack => initInputs_CP_3524_elements(84)); -- 
    -- CP-element group 85:  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_729/if_stmt_833_else_link/$entry
      -- 
    initInputs_CP_3524_elements(85) <= initInputs_CP_3524_elements(82);
    -- CP-element group 86:  transition  input  no-bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_729/if_stmt_833_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_729/if_stmt_833_else_link/else_choice_transition
      -- 
    else_choice_transition_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_833_branch_ack_0, ack => initInputs_CP_3524_elements(86)); -- 
    -- CP-element group 87:  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	200 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_729/xx_x_crit_edge4_xx_x_crit_edge
      -- 
    initInputs_CP_3524_elements(87) <= initInputs_CP_3524_elements(84);
    -- CP-element group 88:  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	187 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_729/xx_x_crit_edge4_bbx_xnph
      -- 
    initInputs_CP_3524_elements(88) <= initInputs_CP_3524_elements(86);
    -- CP-element group 89:  fork  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	12 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	93 
    -- CP-element group 89:  members (10) 
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/$entry
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_update_start_
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_update_start_
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Update/cr
      -- 
    rr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(89), ack => ADD_u16_u16_843_inst_req_0); -- 
    cr_4155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(89), ack => ADD_u16_u16_843_inst_req_1); -- 
    cr_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(89), ack => type_cast_847_inst_req_1); -- 
    initInputs_CP_3524_elements(89) <= initInputs_CP_3524_elements(12);
    -- CP-element group 90:  transition  input  no-bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Sample/ra
      -- 
    ra_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_843_inst_ack_0, ack => initInputs_CP_3524_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  no-bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/ADD_u16_u16_843_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Sample/rr
      -- 
    ca_4156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_843_inst_ack_1, ack => initInputs_CP_3524_elements(91)); -- 
    rr_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(91), ack => type_cast_847_inst_req_0); -- 
    -- CP-element group 92:  transition  input  no-bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Sample/ra
      -- 
    ra_4165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => initInputs_CP_3524_elements(92)); -- 
    -- CP-element group 93:  transition  input  no-bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	89 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	13 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/$exit
      -- CP-element group 93: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_729/assign_stmt_844_to_assign_stmt_848/type_cast_847_Update/ca
      -- 
    ca_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => initInputs_CP_3524_elements(93)); -- 
    -- CP-element group 94:  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_729/do_while_stmt_857/$entry
      -- 
    initInputs_CP_3524_elements(94) <= initInputs_CP_3524_elements(14);
    -- CP-element group 95:  place  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	101 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857__entry__
      -- 
    initInputs_CP_3524_elements(95) <= initInputs_CP_3524_elements(94);
    -- CP-element group 96:  merge  place  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	159 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857__exit__
      -- 
    -- Element group initInputs_CP_3524_elements(96) is bound as output of CP function.
    -- CP-element group 97:  merge  place  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_729/do_while_stmt_857/loop_back
      -- 
    -- Element group initInputs_CP_3524_elements(97) is bound as output of CP function.
    -- CP-element group 98:  branch  place  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	103 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: 	157 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_729/do_while_stmt_857/condition_done
      -- 
    initInputs_CP_3524_elements(98) <= initInputs_CP_3524_elements(103);
    -- CP-element group 99:  branch  place  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	208 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_729/do_while_stmt_857/loop_body_done
      -- 
    initInputs_CP_3524_elements(99) <= initInputs_CP_3524_elements(208);
    -- CP-element group 100:  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	109 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/back_edge_to_loop_body
      -- 
    initInputs_CP_3524_elements(100) <= initInputs_CP_3524_elements(97);
    -- CP-element group 101:  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	95 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	111 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/first_time_through_loop_body
      -- 
    initInputs_CP_3524_elements(101) <= initInputs_CP_3524_elements(95);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	105 
    -- CP-element group 102: 	106 
    -- CP-element group 102: 	128 
    -- CP-element group 102: 	132 
    -- CP-element group 102: 	135 
    -- CP-element group 102: 	140 
    -- CP-element group 102: 	148 
    -- CP-element group 102: 	152 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/$entry
      -- CP-element group 102: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/loop_body_start
      -- 
    -- Element group initInputs_CP_3524_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	106 
    -- CP-element group 103: 	150 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	98 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/condition_evaluated
      -- 
    condition_evaluated_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(103), ack => do_while_stmt_857_branch_req_0); -- 
    initInputs_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 16);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(106) & initInputs_CP_3524_elements(150);
      gj_initInputs_cp_element_group_103 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	108 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/aggregated_phi_sample_req
      -- CP-element group 104: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_sample_start__ps
      -- 
    initInputs_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(105) & initInputs_CP_3524_elements(108);
      gj_initInputs_cp_element_group_104 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  no-bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	146 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	104 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_sample_start_
      -- 
    initInputs_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(107) & initInputs_CP_3524_elements(146);
      gj_initInputs_cp_element_group_105 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  fork  transition  no-bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	102 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: 	129 
    -- CP-element group 106: 	145 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	103 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/aggregated_phi_update_req
      -- CP-element group 106: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_update_start_
      -- CP-element group 106: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_update_start__ps
      -- 
    initInputs_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 16,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(108) & initInputs_CP_3524_elements(129) & initInputs_CP_3524_elements(145);
      gj_initInputs_cp_element_group_106 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	144 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/aggregated_phi_sample_ack
      -- CP-element group 107: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_sample_completed__ps
      -- 
    -- Element group initInputs_CP_3524_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	127 
    -- CP-element group 108: 	143 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/aggregated_phi_update_ack
      -- CP-element group 108: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_update_completed__ps
      -- 
    -- Element group initInputs_CP_3524_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	100 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_loopback_trigger
      -- 
    initInputs_CP_3524_elements(109) <= initInputs_CP_3524_elements(100);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	115 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_loopback_sample_req
      -- 
    phi_stmt_859_loopback_sample_req_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_859_loopback_sample_req_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(110), ack => phi_stmt_859_req_0); -- 
    -- Element group initInputs_CP_3524_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	101 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_entry_trigger
      -- 
    initInputs_CP_3524_elements(111) <= initInputs_CP_3524_elements(101);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_entry_sample_req
      -- 
    phi_stmt_859_entry_sample_req_4202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_859_entry_sample_req_4202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(112), ack => phi_stmt_859_req_1); -- 
    -- Element group initInputs_CP_3524_elements(112) is bound as output of CP function.
    -- CP-element group 113:  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_merged_reqs
      -- 
    -- Element group initInputs_CP_3524_elements(113) is bound as output of CP function.
    -- CP-element group 114:  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_entry_sample_req__merge_in
      -- 
    initInputs_CP_3524_elements(114) <= initInputs_CP_3524_elements(112);
    -- CP-element group 115:  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	110 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_loopback_sample_req__merge_in
      -- 
    initInputs_CP_3524_elements(115) <= initInputs_CP_3524_elements(110);
    -- CP-element group 116:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	208 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_phi_mux_ack
      -- 
    phi_stmt_859_phi_mux_ack_4207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_859_ack_0, ack => initInputs_CP_3524_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_sample_start__ps
      -- 
    -- Element group initInputs_CP_3524_elements(117) is bound as output of CP function.
    -- CP-element group 118:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_update_start__ps
      -- 
    -- Element group initInputs_CP_3524_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Sample/rr
      -- 
    rr_4220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(119), ack => type_cast_862_inst_req_0); -- 
    initInputs_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(117) & initInputs_CP_3524_elements(121);
      gj_initInputs_cp_element_group_119 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_update_start_
      -- CP-element group 120: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Update/cr
      -- 
    cr_4225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(120), ack => type_cast_862_inst_req_1); -- 
    initInputs_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(118) & initInputs_CP_3524_elements(122);
      gj_initInputs_cp_element_group_120 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Sample/ra
      -- 
    ra_4221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_0, ack => initInputs_CP_3524_elements(121)); -- 
    -- CP-element group 122:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_update_completed__ps
      -- CP-element group 122: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/type_cast_862_Update/ca
      -- 
    ca_4226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_1, ack => initInputs_CP_3524_elements(122)); -- 
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_sample_start__ps
      -- CP-element group 123: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Sample/req
      -- 
    req_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(123), ack => indvar_at_entry_851_863_buf_req_0); -- 
    -- Element group initInputs_CP_3524_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_update_start__ps
      -- CP-element group 124: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_update_start_
      -- CP-element group 124: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Update/req
      -- 
    req_4243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(124), ack => indvar_at_entry_851_863_buf_req_1); -- 
    -- Element group initInputs_CP_3524_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Sample/ack
      -- 
    ack_4239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => indvar_at_entry_851_863_buf_ack_0, ack => initInputs_CP_3524_elements(125)); -- 
    -- CP-element group 126:  join  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_update_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/R_indvar_at_entry_863_Update/ack
      -- 
    ack_4244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => indvar_at_entry_851_863_buf_ack_1, ack => initInputs_CP_3524_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	108 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Sample/rr
      -- 
    rr_4253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(127), ack => ADD_u64_u64_869_inst_req_0); -- 
    initInputs_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(108) & initInputs_CP_3524_elements(129);
      gj_initInputs_cp_element_group_127 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	102 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_update_start_
      -- CP-element group 128: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Update/cr
      -- 
    cr_4258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(128), ack => ADD_u64_u64_869_inst_req_1); -- 
    initInputs_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(130);
      gj_initInputs_cp_element_group_128 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	106 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Sample/ra
      -- 
    ra_4254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_869_inst_ack_0, ack => initInputs_CP_3524_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (24) 
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_869_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_root_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_offset_calculated
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_resized_0
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_scaled_0
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_computed_0
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_resize_0/$entry
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_resize_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_resize_0/index_resize_req
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_resize_0/index_resize_ack
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_scale_0/$entry
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_scale_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_scale_0/scale_rename_req
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_index_scale_0/scale_rename_ack
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_final_index_sum_regn/$entry
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_final_index_sum_regn/$exit
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_final_index_sum_regn/req
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_final_index_sum_regn/ack
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_base_plus_offset/$entry
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_base_plus_offset/$exit
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_base_plus_offset/sum_rename_req
      -- CP-element group 130: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/array_obj_ref_873_base_plus_offset/sum_rename_ack
      -- 
    ca_4259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_869_inst_ack_1, ack => initInputs_CP_3524_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_request/$entry
      -- CP-element group 131: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_request/req
      -- 
    req_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(131), ack => addr_of_874_final_reg_req_0); -- 
    initInputs_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(130) & initInputs_CP_3524_elements(133);
      gj_initInputs_cp_element_group_131 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	102 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	141 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_update_start_
      -- CP-element group 132: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_complete/$entry
      -- CP-element group 132: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_complete/req
      -- 
    req_4297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(132), ack => addr_of_874_final_reg_req_1); -- 
    initInputs_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(134) & initInputs_CP_3524_elements(141);
      gj_initInputs_cp_element_group_132 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	208 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_request/$exit
      -- CP-element group 133: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_request/ack
      -- 
    ack_4293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_874_final_reg_ack_0, ack => initInputs_CP_3524_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	139 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (19) 
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/addr_of_874_complete/ack
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_word_addrgen/root_register_ack
      -- 
    ack_4298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_874_final_reg_ack_1, ack => initInputs_CP_3524_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	102 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Sample/rr
      -- 
    rr_4306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(135), ack => RPIPE_matrix_in_877_inst_req_0); -- 
    initInputs_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(137);
      gj_initInputs_cp_element_group_135 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: 	141 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_update_start_
      -- CP-element group 136: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Update/cr
      -- 
    cr_4311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(136), ack => RPIPE_matrix_in_877_inst_req_1); -- 
    initInputs_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(137) & initInputs_CP_3524_elements(138) & initInputs_CP_3524_elements(141);
      gj_initInputs_cp_element_group_136 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Sample/ra
      -- 
    ra_4307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_877_inst_ack_0, ack => initInputs_CP_3524_elements(137)); -- 
    -- CP-element group 138:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/RPIPE_matrix_in_877_Update/ca
      -- 
    ca_4312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_matrix_in_877_inst_ack_1, ack => initInputs_CP_3524_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	134 
    -- CP-element group 139: 	138 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/ptr_deref_880_Split/$entry
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/ptr_deref_880_Split/$exit
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/ptr_deref_880_Split/split_req
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/ptr_deref_880_Split/split_ack
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/$entry
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/word_0/$entry
      -- CP-element group 139: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/word_0/rr
      -- 
    rr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(139), ack => ptr_deref_880_store_0_req_0); -- 
    initInputs_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 16,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(134) & initInputs_CP_3524_elements(138) & initInputs_CP_3524_elements(141);
      gj_initInputs_cp_element_group_139 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	102 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (5) 
      -- CP-element group 140: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_update_start_
      -- CP-element group 140: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/$entry
      -- CP-element group 140: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/word_0/$entry
      -- CP-element group 140: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/word_0/cr
      -- 
    cr_4361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(140), ack => ptr_deref_880_store_0_req_1); -- 
    initInputs_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(142);
      gj_initInputs_cp_element_group_140 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	132 
    -- CP-element group 141: 	136 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (5) 
      -- CP-element group 141: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/$exit
      -- CP-element group 141: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/word_0/$exit
      -- CP-element group 141: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Sample/word_access_start/word_0/ra
      -- 
    ra_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_0, ack => initInputs_CP_3524_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	208 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/word_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ptr_deref_880_Update/word_access_complete/word_0/ca
      -- 
    ca_4362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_1, ack => initInputs_CP_3524_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	108 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Sample/rr
      -- 
    rr_4370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(143), ack => ADD_u64_u64_887_inst_req_0); -- 
    initInputs_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(108) & initInputs_CP_3524_elements(145);
      gj_initInputs_cp_element_group_143 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	107 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: 	149 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_update_start_
      -- CP-element group 144: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Update/cr
      -- 
    cr_4375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(144), ack => ADD_u64_u64_887_inst_req_1); -- 
    initInputs_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(107) & initInputs_CP_3524_elements(146) & initInputs_CP_3524_elements(149);
      gj_initInputs_cp_element_group_144 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	106 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Sample/ra
      -- 
    ra_4371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_887_inst_ack_0, ack => initInputs_CP_3524_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	105 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/ADD_u64_u64_887_Update/ca
      -- 
    ca_4376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_887_inst_ack_1, ack => initInputs_CP_3524_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Sample/rr
      -- 
    rr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(147), ack => EQ_u64_u1_892_inst_req_0); -- 
    initInputs_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(146) & initInputs_CP_3524_elements(149);
      gj_initInputs_cp_element_group_147 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	102 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_update_start_
      -- CP-element group 148: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Update/cr
      -- 
    cr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(148), ack => EQ_u64_u1_892_inst_req_1); -- 
    initInputs_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(150) & initInputs_CP_3524_elements(153);
      gj_initInputs_cp_element_group_148 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	144 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Sample/ra
      -- 
    ra_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_892_inst_ack_0, ack => initInputs_CP_3524_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	103 
    -- CP-element group 150: 	151 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/EQ_u64_u1_892_Update/ca
      -- 
    ca_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_892_inst_ack_1, ack => initInputs_CP_3524_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Sample/req
      -- 
    req_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(151), ack => W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_0); -- 
    initInputs_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(150) & initInputs_CP_3524_elements(153);
      gj_initInputs_cp_element_group_151 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	102 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_update_start_
      -- CP-element group 152: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Update/req
      -- 
    req_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(152), ack => W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_1); -- 
    initInputs_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(102) & initInputs_CP_3524_elements(154);
      gj_initInputs_cp_element_group_152 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Sample/ack
      -- 
    ack_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_0, ack => initInputs_CP_3524_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	208 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/assign_stmt_896_Update/ack
      -- 
    ack_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_1, ack => initInputs_CP_3524_elements(154)); -- 
    -- CP-element group 155:  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	98 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_729/do_while_stmt_857/loop_exit/$entry
      -- 
    initInputs_CP_3524_elements(155) <= initInputs_CP_3524_elements(98);
    -- CP-element group 156:  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_729/do_while_stmt_857/loop_exit/$exit
      -- CP-element group 156: 	 branch_block_stmt_729/do_while_stmt_857/loop_exit/ack
      -- 
    ack_4408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_857_branch_ack_0, ack => initInputs_CP_3524_elements(156)); -- 
    -- CP-element group 157:  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	98 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_729/do_while_stmt_857/loop_taken/$entry
      -- 
    initInputs_CP_3524_elements(157) <= initInputs_CP_3524_elements(98);
    -- CP-element group 158:  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_729/do_while_stmt_857/loop_taken/$exit
      -- CP-element group 158: 	 branch_block_stmt_729/do_while_stmt_857/loop_taken/ack
      -- 
    ack_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_857_branch_ack_1, ack => initInputs_CP_3524_elements(158)); -- 
    -- CP-element group 159:  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	96 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	15 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_729/do_while_stmt_857/$exit
      -- 
    initInputs_CP_3524_elements(159) <= initInputs_CP_3524_elements(96);
    -- CP-element group 160:  transition  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	15 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_729/if_stmt_900_dead_link/$entry
      -- 
    initInputs_CP_3524_elements(160) <= initInputs_CP_3524_elements(15);
    -- CP-element group 161:  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	15 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_729/if_stmt_900_eval_test/$entry
      -- CP-element group 161: 	 branch_block_stmt_729/if_stmt_900_eval_test/$exit
      -- CP-element group 161: 	 branch_block_stmt_729/if_stmt_900_eval_test/branch_req
      -- 
    branch_req_4421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(161), ack => if_stmt_900_branch_req_0); -- 
    initInputs_CP_3524_elements(161) <= initInputs_CP_3524_elements(15);
    -- CP-element group 162:  branch  place  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	165 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_729/R_bb_4_xx_x_crit_edgex_xloopexit_taken_901_place
      -- 
    initInputs_CP_3524_elements(162) <= initInputs_CP_3524_elements(161);
    -- CP-element group 163:  transition  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_729/if_stmt_900_if_link/$entry
      -- 
    initInputs_CP_3524_elements(163) <= initInputs_CP_3524_elements(162);
    -- CP-element group 164:  transition  input  no-bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	167 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_729/if_stmt_900_if_link/$exit
      -- CP-element group 164: 	 branch_block_stmt_729/if_stmt_900_if_link/if_choice_transition
      -- 
    if_choice_transition_4426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_900_branch_ack_1, ack => initInputs_CP_3524_elements(164)); -- 
    -- CP-element group 165:  transition  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_729/if_stmt_900_else_link/$entry
      -- 
    initInputs_CP_3524_elements(165) <= initInputs_CP_3524_elements(162);
    -- CP-element group 166:  transition  input  no-bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	16 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_729/if_stmt_900_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_729/if_stmt_900_else_link/else_choice_transition
      -- 
    else_choice_transition_4430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_900_branch_ack_0, ack => initInputs_CP_3524_elements(166)); -- 
    -- CP-element group 167:  place  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	164 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	197 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_729/bb_4_xx_x_crit_edgex_xloopexit
      -- 
    initInputs_CP_3524_elements(167) <= initInputs_CP_3524_elements(164);
    -- CP-element group 168:  transition  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	18 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_729/assign_stmt_909/$entry
      -- CP-element group 168: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Sample/rr
      -- 
    rr_4442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(168), ack => RPIPE_rate_in_908_inst_req_0); -- 
    initInputs_CP_3524_elements(168) <= initInputs_CP_3524_elements(18);
    -- CP-element group 169:  transition  input  output  no-bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_update_start_
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Sample/ra
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Update/cr
      -- 
    ra_4443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rate_in_908_inst_ack_0, ack => initInputs_CP_3524_elements(169)); -- 
    cr_4447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(169), ack => RPIPE_rate_in_908_inst_req_1); -- 
    -- CP-element group 170:  transition  input  no-bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	19 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_729/assign_stmt_909/$exit
      -- CP-element group 170: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_729/assign_stmt_909/RPIPE_rate_in_908_Update/ca
      -- 
    ca_4448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rate_in_908_inst_ack_1, ack => initInputs_CP_3524_elements(170)); -- 
    -- CP-element group 171:  fork  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	19 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (17) 
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_update_start_
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_word_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/STORE_rate_910_Split/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/STORE_rate_910_Split/$exit
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/STORE_rate_910_Split/split_req
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/STORE_rate_910_Split/split_ack
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/word_0/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/word_0/rr
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/word_0/$entry
      -- CP-element group 171: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/word_0/cr
      -- 
    cr_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(171), ack => STORE_rate_910_store_0_req_1); -- 
    rr_4472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(171), ack => STORE_rate_910_store_0_req_0); -- 
    initInputs_CP_3524_elements(171) <= initInputs_CP_3524_elements(19);
    -- CP-element group 172:  transition  input  no-bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (5) 
      -- CP-element group 172: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/$exit
      -- CP-element group 172: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/word_0/$exit
      -- CP-element group 172: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Sample/word_access_start/word_0/ra
      -- 
    ra_4473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_rate_910_store_0_ack_0, ack => initInputs_CP_3524_elements(172)); -- 
    -- CP-element group 173:  transition  input  no-bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	20 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/$exit
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/word_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_729/assign_stmt_912/STORE_rate_910_Update/word_access_complete/word_0/ca
      -- 
    ca_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_rate_910_store_0_ack_1, ack => initInputs_CP_3524_elements(173)); -- 
    -- CP-element group 174:  fork  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	57 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Update/cr
      -- 
    rr_4503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(174), ack => type_cast_750_inst_req_0); -- 
    cr_4508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(174), ack => type_cast_750_inst_req_1); -- 
    initInputs_CP_3524_elements(174) <= initInputs_CP_3524_elements(57);
    -- CP-element group 175:  transition  input  no-bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Sample/ra
      -- 
    ra_4504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => initInputs_CP_3524_elements(175)); -- 
    -- CP-element group 176:  transition  input  no-bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/Update/ca
      -- 
    ca_4509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => initInputs_CP_3524_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	181 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/$exit
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/$exit
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/$exit
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/$exit
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_750/SplitProtocol/$exit
      -- CP-element group 177: 	 branch_block_stmt_729/bb_1_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_req
      -- 
    phi_stmt_744_req_4510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_744_req_4510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(177), ack => phi_stmt_744_req_1); -- 
    initInputs_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(175) & initInputs_CP_3524_elements(176);
      gj_initInputs_cp_element_group_177 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	5 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/$entry
      -- CP-element group 178: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/$entry
      -- CP-element group 178: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/$entry
      -- 
    initInputs_CP_3524_elements(178) <= initInputs_CP_3524_elements(5);
    -- CP-element group 179:  transition  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/type_cast_748_konst_delay_trans
      -- 
    -- Element group initInputs_CP_3524_elements(179) is a control-delay.
    cp_element_179_delay: control_delay_element  generic map(name => " 179_delay", delay_value => 1)  port map(req => initInputs_CP_3524_elements(178), ack => initInputs_CP_3524_elements(179), clk => clk, reset =>reset);
    -- CP-element group 180:  transition  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (4) 
      -- CP-element group 180: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/$exit
      -- CP-element group 180: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/$exit
      -- CP-element group 180: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_sources/$exit
      -- CP-element group 180: 	 branch_block_stmt_729/bbx_xnph3_bb_1_PhiReq/phi_stmt_744/phi_stmt_744_req
      -- 
    phi_stmt_744_req_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_744_req_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(180), ack => phi_stmt_744_req_0); -- 
    initInputs_CP_3524_elements(180) <= initInputs_CP_3524_elements(179);
    -- CP-element group 181:  merge  place  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	177 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_729/merge_stmt_743_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(181) <= OrReduce(initInputs_CP_3524_elements(177) & initInputs_CP_3524_elements(180));
    -- CP-element group 182:  transition  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_729/merge_stmt_743_PhiAck/$entry
      -- 
    initInputs_CP_3524_elements(182) <= initInputs_CP_3524_elements(181);
    -- CP-element group 183:  transition  input  no-bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	6 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_729/merge_stmt_743_PhiAck/$exit
      -- CP-element group 183: 	 branch_block_stmt_729/merge_stmt_743_PhiAck/phi_stmt_744_ack
      -- 
    phi_stmt_744_ack_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_744_ack_0, ack => initInputs_CP_3524_elements(183)); -- 
    -- CP-element group 184:  transition  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	56 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_729/bb_1_xx_x_crit_edge4_PhiReq/$entry
      -- CP-element group 184: 	 branch_block_stmt_729/bb_1_xx_x_crit_edge4_PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(184) <= initInputs_CP_3524_elements(56);
    -- CP-element group 185:  place  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_729/merge_stmt_782_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(185) <= initInputs_CP_3524_elements(184);
    -- CP-element group 186:  transition  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	10 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_729/merge_stmt_782_PhiAck/$entry
      -- CP-element group 186: 	 branch_block_stmt_729/merge_stmt_782_PhiAck/$exit
      -- CP-element group 186: 	 branch_block_stmt_729/merge_stmt_782_PhiAck/dummy
      -- 
    initInputs_CP_3524_elements(186) <= initInputs_CP_3524_elements(185);
    -- CP-element group 187:  transition  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	88 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_729/xx_x_crit_edge4_bbx_xnph_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_729/xx_x_crit_edge4_bbx_xnph_PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(187) <= initInputs_CP_3524_elements(88);
    -- CP-element group 188:  place  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_729/merge_stmt_839_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(188) <= initInputs_CP_3524_elements(187);
    -- CP-element group 189:  transition  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	12 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_729/merge_stmt_839_PhiAck/$entry
      -- CP-element group 189: 	 branch_block_stmt_729/merge_stmt_839_PhiAck/$exit
      -- CP-element group 189: 	 branch_block_stmt_729/merge_stmt_839_PhiAck/dummy
      -- 
    initInputs_CP_3524_elements(189) <= initInputs_CP_3524_elements(188);
    -- CP-element group 190:  transition  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	13 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/$entry
      -- CP-element group 190: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/$entry
      -- CP-element group 190: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/phi_stmt_851_sources/$entry
      -- 
    initInputs_CP_3524_elements(190) <= initInputs_CP_3524_elements(13);
    -- CP-element group 191:  transition  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/phi_stmt_851_sources/type_cast_855_konst_delay_trans
      -- 
    -- Element group initInputs_CP_3524_elements(191) is a control-delay.
    cp_element_191_delay: control_delay_element  generic map(name => " 191_delay", delay_value => 1)  port map(req => initInputs_CP_3524_elements(190), ack => initInputs_CP_3524_elements(191), clk => clk, reset =>reset);
    -- CP-element group 192:  transition  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (4) 
      -- CP-element group 192: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/$exit
      -- CP-element group 192: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/$exit
      -- CP-element group 192: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/phi_stmt_851_sources/$exit
      -- CP-element group 192: 	 branch_block_stmt_729/bbx_xnph_bb_4_PhiReq/phi_stmt_851/phi_stmt_851_req
      -- 
    phi_stmt_851_req_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_851_req_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initInputs_CP_3524_elements(192), ack => phi_stmt_851_req_0); -- 
    initInputs_CP_3524_elements(192) <= initInputs_CP_3524_elements(191);
    -- CP-element group 193:  place  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_729/merge_stmt_850_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(193) <= initInputs_CP_3524_elements(192);
    -- CP-element group 194:  transition  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_729/merge_stmt_850_PhiAck/$entry
      -- 
    initInputs_CP_3524_elements(194) <= initInputs_CP_3524_elements(193);
    -- CP-element group 195:  transition  input  no-bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	14 
    -- CP-element group 195:  members (2) 
      -- CP-element group 195: 	 branch_block_stmt_729/merge_stmt_850_PhiAck/$exit
      -- CP-element group 195: 	 branch_block_stmt_729/merge_stmt_850_PhiAck/phi_stmt_851_ack
      -- 
    phi_stmt_851_ack_4566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_851_ack_0, ack => initInputs_CP_3524_elements(195)); -- 
    -- CP-element group 196:  transition  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	16 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_729/merge_stmt_904_dead_link/$entry
      -- 
    initInputs_CP_3524_elements(196) <= initInputs_CP_3524_elements(16);
    -- CP-element group 197:  transition  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	167 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_729/bb_4_xx_x_crit_edgex_xloopexit_PhiReq/$entry
      -- CP-element group 197: 	 branch_block_stmt_729/bb_4_xx_x_crit_edgex_xloopexit_PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(197) <= initInputs_CP_3524_elements(167);
    -- CP-element group 198:  place  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_729/merge_stmt_904_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(198) <= initInputs_CP_3524_elements(197);
    -- CP-element group 199:  transition  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	17 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_729/merge_stmt_904_PhiAck/$entry
      -- CP-element group 199: 	 branch_block_stmt_729/merge_stmt_904_PhiAck/$exit
      -- CP-element group 199: 	 branch_block_stmt_729/merge_stmt_904_PhiAck/dummy
      -- 
    initInputs_CP_3524_elements(199) <= initInputs_CP_3524_elements(198);
    -- CP-element group 200:  transition  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	87 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_729/xx_x_crit_edge4_xx_x_crit_edge_PhiReq/$entry
      -- CP-element group 200: 	 branch_block_stmt_729/xx_x_crit_edge4_xx_x_crit_edge_PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(200) <= initInputs_CP_3524_elements(87);
    -- CP-element group 201:  transition  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	17 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_729/xx_x_crit_edgex_xloopexit_xx_x_crit_edge_PhiReq/$entry
      -- CP-element group 201: 	 branch_block_stmt_729/xx_x_crit_edgex_xloopexit_xx_x_crit_edge_PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(201) <= initInputs_CP_3524_elements(17);
    -- CP-element group 202:  merge  place  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_729/merge_stmt_906_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(202) <= OrReduce(initInputs_CP_3524_elements(200) & initInputs_CP_3524_elements(201));
    -- CP-element group 203:  transition  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	18 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_729/merge_stmt_906_PhiAck/$entry
      -- CP-element group 203: 	 branch_block_stmt_729/merge_stmt_906_PhiAck/$exit
      -- CP-element group 203: 	 branch_block_stmt_729/merge_stmt_906_PhiAck/dummy
      -- 
    initInputs_CP_3524_elements(203) <= initInputs_CP_3524_elements(202);
    -- CP-element group 204:  transition  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	20 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (2) 
      -- CP-element group 204: 	 branch_block_stmt_729/return___PhiReq/$entry
      -- CP-element group 204: 	 branch_block_stmt_729/return___PhiReq/$exit
      -- 
    initInputs_CP_3524_elements(204) <= initInputs_CP_3524_elements(20);
    -- CP-element group 205:  place  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_729/merge_stmt_914_PhiReqMerge
      -- 
    initInputs_CP_3524_elements(205) <= initInputs_CP_3524_elements(204);
    -- CP-element group 206:  transition  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	21 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_729/merge_stmt_914_PhiAck/$entry
      -- CP-element group 206: 	 branch_block_stmt_729/merge_stmt_914_PhiAck/$exit
      -- CP-element group 206: 	 branch_block_stmt_729/merge_stmt_914_PhiAck/dummy
      -- 
    initInputs_CP_3524_elements(206) <= initInputs_CP_3524_elements(205);
    -- CP-element group 207:  transition  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	21 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (2) 
      -- CP-element group 207: 	 $exit
      -- CP-element group 207: 	 branch_block_stmt_729/$exit
      -- 
    initInputs_CP_3524_elements(207) <= initInputs_CP_3524_elements(21);
    -- CP-element group 208:  join  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	116 
    -- CP-element group 208: 	133 
    -- CP-element group 208: 	142 
    -- CP-element group 208: 	154 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	99 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/$exit
      -- CP-element group 208: 	 branch_block_stmt_729/do_while_stmt_857/do_while_stmt_857_loop_body/phi_stmt_859_phi_mux_ack_ps
      -- 
    initInputs_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 16,1 => 16,2 => 16,3 => 16);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "initInputs_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= initInputs_CP_3524_elements(116) & initInputs_CP_3524_elements(133) & initInputs_CP_3524_elements(142) & initInputs_CP_3524_elements(154);
      gj_initInputs_cp_element_group_208 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initInputs_CP_3524_elements(208), clk => clk, reset => reset); --
    end block;
    initInputs_do_while_stmt_857_terminator_4413: loop_terminator -- 
      generic map (name => " initInputs_do_while_stmt_857_terminator_4413", max_iterations_in_flight =>16) 
      port map(loop_body_exit => initInputs_CP_3524_elements(99),loop_continue => initInputs_CP_3524_elements(158),loop_terminate => initInputs_CP_3524_elements(156),loop_back => initInputs_CP_3524_elements(97),loop_exit => initInputs_CP_3524_elements(96),clk => clk, reset => reset); -- 
    phi_stmt_859_phi_seq_4245_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initInputs_CP_3524_elements(109);
      initInputs_CP_3524_elements(117)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initInputs_CP_3524_elements(121);
      initInputs_CP_3524_elements(118)<= src_update_reqs(0);
      src_update_acks(0)  <= initInputs_CP_3524_elements(122);
      initInputs_CP_3524_elements(110) <= phi_mux_reqs(0);
      triggers(1)  <= initInputs_CP_3524_elements(111);
      initInputs_CP_3524_elements(123)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initInputs_CP_3524_elements(125);
      initInputs_CP_3524_elements(124)<= src_update_reqs(1);
      src_update_acks(1)  <= initInputs_CP_3524_elements(126);
      initInputs_CP_3524_elements(112) <= phi_mux_reqs(1);
      phi_stmt_859_phi_seq_4245 : phi_sequencer_v2-- 
        generic map (place_capacity => 16, ntriggers => 2, name => "phi_stmt_859_phi_seq_4245") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initInputs_CP_3524_elements(104), 
          phi_sample_ack => initInputs_CP_3524_elements(107), 
          phi_update_req => initInputs_CP_3524_elements(106), 
          phi_update_ack => initInputs_CP_3524_elements(108), 
          phi_mux_ack => initInputs_CP_3524_elements(116), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4186_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= initInputs_CP_3524_elements(100);
        preds(1)  <= initInputs_CP_3524_elements(101);
        entry_tmerge_4186 : transition_merge -- 
          generic map(name => " entry_tmerge_4186")
          port map (preds => preds, symbol_out => initInputs_CP_3524_elements(102));
          -- 
    end block;
    phi_stmt_859_req_merge_4206_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= initInputs_CP_3524_elements(114);
        preds(1)  <= initInputs_CP_3524_elements(115);
        phi_stmt_859_req_merge_4206 : transition_merge -- 
          generic map(name => " phi_stmt_859_req_merge_4206")
          port map (preds => preds, symbol_out => initInputs_CP_3524_elements(113));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_899_wire : std_logic_vector(0 downto 0);
    signal R_indvar7_753_resized : std_logic_vector(9 downto 0);
    signal R_indvar7_753_scaled : std_logic_vector(9 downto 0);
    signal R_tmp3_872_resized : std_logic_vector(9 downto 0);
    signal R_tmp3_872_scaled : std_logic_vector(9 downto 0);
    signal STORE_ebbyNo_739_data_0 : std_logic_vector(31 downto 0);
    signal STORE_ebbyNo_739_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_maxNitr_733_data_0 : std_logic_vector(15 downto 0);
    signal STORE_maxNitr_733_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ncol_ind_819_data_0 : std_logic_vector(15 downto 0);
    signal STORE_ncol_ind_819_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ncols_806_data_0 : std_logic_vector(15 downto 0);
    signal STORE_ncols_806_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_nrows_793_data_0 : std_logic_vector(15 downto 0);
    signal STORE_nrows_793_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_rate_910_data_0 : std_logic_vector(31 downto 0);
    signal STORE_rate_910_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_754_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_754_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_754_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_754_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_873_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_873_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_873_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_873_root_address : std_logic_vector(9 downto 0);
    signal bb_4_xx_x_crit_edgex_xloopexit_taken_896 : std_logic_vector(0 downto 0);
    signal exitcond2_893 : std_logic_vector(0 downto 0);
    signal exitcond_775 : std_logic_vector(0 downto 0);
    signal iNsTr_11_788 : std_logic_vector(31 downto 0);
    signal iNsTr_12_792 : std_logic_vector(15 downto 0);
    signal iNsTr_14_801 : std_logic_vector(31 downto 0);
    signal iNsTr_15_805 : std_logic_vector(15 downto 0);
    signal iNsTr_17_814 : std_logic_vector(31 downto 0);
    signal iNsTr_18_818 : std_logic_vector(15 downto 0);
    signal iNsTr_1_732 : std_logic_vector(15 downto 0);
    signal iNsTr_20_827 : std_logic_vector(15 downto 0);
    signal iNsTr_21_832 : std_logic_vector(0 downto 0);
    signal iNsTr_24_909 : std_logic_vector(31 downto 0);
    signal iNsTr_30_878 : std_logic_vector(15 downto 0);
    signal iNsTr_4_738 : std_logic_vector(31 downto 0);
    signal iNsTr_8_759 : std_logic_vector(15 downto 0);
    signal indvar7_744 : std_logic_vector(63 downto 0);
    signal indvar_859 : std_logic_vector(63 downto 0);
    signal indvar_at_entry_851 : std_logic_vector(63 downto 0);
    signal indvar_at_entry_851_863_buffered : std_logic_vector(63 downto 0);
    signal indvarx_xnext8_769 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_888 : std_logic_vector(63 downto 0);
    signal ptr_deref_761_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_761_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_761_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_761_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_761_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_761_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_791_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_791_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_791_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_791_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_791_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_804_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_804_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_804_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_804_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_804_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_817_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_817_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_817_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_817_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_817_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_880_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_880_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_880_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_880_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_880_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_880_word_offset_0 : std_logic_vector(9 downto 0);
    signal scevgep10_756 : std_logic_vector(31 downto 0);
    signal scevgep_875 : std_logic_vector(31 downto 0);
    signal tmp1_848 : std_logic_vector(63 downto 0);
    signal tmp3_870 : std_logic_vector(63 downto 0);
    signal tmp_844 : std_logic_vector(15 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_750_wire : std_logic_vector(63 downto 0);
    signal type_cast_767_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_855_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_862_wire : std_logic_vector(63 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_ebbyNo_739_word_address_0 <= "0";
    STORE_maxNitr_733_word_address_0 <= "0";
    STORE_ncol_ind_819_word_address_0 <= "0";
    STORE_ncols_806_word_address_0 <= "0";
    STORE_nrows_793_word_address_0 <= "0";
    STORE_rate_910_word_address_0 <= "0";
    array_obj_ref_754_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_754_resized_base_address <= "0000000000";
    array_obj_ref_873_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_873_resized_base_address <= "0000000000";
    iNsTr_11_788 <= "00000000000000000000000000000000";
    iNsTr_14_801 <= "00000000000000000000000000000001";
    iNsTr_17_814 <= "00000000000000000000000000000010";
    ptr_deref_761_word_offset_0 <= "0000000000";
    ptr_deref_791_word_offset_0 <= "0000000000";
    ptr_deref_804_word_offset_0 <= "0000000000";
    ptr_deref_817_word_offset_0 <= "0000000000";
    ptr_deref_880_word_offset_0 <= "0000000000";
    type_cast_748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_767_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_824_wire_constant <= "0000000000000000";
    type_cast_855_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_868_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_886_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_744: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_748_wire_constant & type_cast_750_wire;
      req <= phi_stmt_744_req_0 & phi_stmt_744_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_744",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_744_ack_0,
          idata => idata,
          odata => indvar7_744,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_744
    phi_stmt_851: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_855_wire_constant;
      req(0) <= phi_stmt_851_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_851",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_851_ack_0,
          idata => idata,
          odata => indvar_at_entry_851,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_851
    phi_stmt_859: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_862_wire & indvar_at_entry_851_863_buffered;
      req <= phi_stmt_859_req_0 & phi_stmt_859_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_859",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_859_ack_0,
          idata => idata,
          odata => indvar_859,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_859
    W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_0;
      W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_0<= wack(0);
      rreq(0) <= W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_req_1;
      W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst_ack_1<= rack(0);
      W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst : InterlockBuffer generic map ( -- 
        name => "W_bb_4_xx_x_crit_edgex_xloopexit_taken_894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exitcond2_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bb_4_xx_x_crit_edgex_xloopexit_taken_896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_755_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_755_final_reg_req_0;
      addr_of_755_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_755_final_reg_req_1;
      addr_of_755_final_reg_ack_1<= rack(0);
      addr_of_755_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_755_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_754_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep10_756,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_874_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_874_final_reg_req_0;
      addr_of_874_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_874_final_reg_req_1;
      addr_of_874_final_reg_ack_1<= rack(0);
      addr_of_874_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_874_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_873_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep_875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    indvar_at_entry_851_863_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= indvar_at_entry_851_863_buf_req_0;
      indvar_at_entry_851_863_buf_ack_0<= wack(0);
      rreq(0) <= indvar_at_entry_851_863_buf_req_1;
      indvar_at_entry_851_863_buf_ack_1<= rack(0);
      indvar_at_entry_851_863_buf : InterlockBuffer generic map ( -- 
        name => "indvar_at_entry_851_863_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_at_entry_851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => indvar_at_entry_851_863_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext8_769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_750_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_862_inst_req_0;
      type_cast_862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_862_inst_req_1;
      type_cast_862_inst_ack_1<= rack(0);
      type_cast_862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_888,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_862_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_ebbyNo_739_gather_scatter
    process(iNsTr_4_738) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_738;
      ov(31 downto 0) := iv;
      STORE_ebbyNo_739_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_maxNitr_733_gather_scatter
    process(iNsTr_1_732) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_732;
      ov(15 downto 0) := iv;
      STORE_maxNitr_733_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_ncol_ind_819_gather_scatter
    process(iNsTr_18_818) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_818;
      ov(15 downto 0) := iv;
      STORE_ncol_ind_819_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_ncols_806_gather_scatter
    process(iNsTr_15_805) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_805;
      ov(15 downto 0) := iv;
      STORE_ncols_806_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_nrows_793_gather_scatter
    process(iNsTr_12_792) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_12_792;
      ov(15 downto 0) := iv;
      STORE_nrows_793_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_rate_910_gather_scatter
    process(iNsTr_24_909) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_24_909;
      ov(31 downto 0) := iv;
      STORE_rate_910_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_754_index_0_rename
    process(R_indvar7_753_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar7_753_resized;
      ov(9 downto 0) := iv;
      R_indvar7_753_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_754_index_0_resize
    process(indvar7_744) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar7_744;
      ov := iv(9 downto 0);
      R_indvar7_753_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_754_index_offset
    process(R_indvar7_753_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar7_753_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_754_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_754_root_address_inst
    process(array_obj_ref_754_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_754_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_754_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_873_index_0_rename
    process(R_tmp3_872_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp3_872_resized;
      ov(9 downto 0) := iv;
      R_tmp3_872_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_873_index_0_resize
    process(tmp3_870) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp3_870;
      ov := iv(9 downto 0);
      R_tmp3_872_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_873_index_offset
    process(R_tmp3_872_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp3_872_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_873_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_873_root_address_inst
    process(array_obj_ref_873_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_873_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_873_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_761_addr_0
    process(ptr_deref_761_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_761_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_761_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_761_base_resize
    process(scevgep10_756) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep10_756;
      ov := iv(9 downto 0);
      ptr_deref_761_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_761_gather_scatter
    process(iNsTr_8_759) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_759;
      ov(15 downto 0) := iv;
      ptr_deref_761_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_761_root_address_inst
    process(ptr_deref_761_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_761_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_761_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_791_addr_0
    process(ptr_deref_791_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_791_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_791_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_791_base_resize
    process(iNsTr_11_788) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_11_788;
      ov := iv(9 downto 0);
      ptr_deref_791_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_791_gather_scatter
    process(ptr_deref_791_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_791_data_0;
      ov(15 downto 0) := iv;
      iNsTr_12_792 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_791_root_address_inst
    process(ptr_deref_791_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_791_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_791_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_addr_0
    process(ptr_deref_804_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_804_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_base_resize
    process(iNsTr_14_801) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_14_801;
      ov := iv(9 downto 0);
      ptr_deref_804_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_gather_scatter
    process(ptr_deref_804_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_data_0;
      ov(15 downto 0) := iv;
      iNsTr_15_805 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_804_root_address_inst
    process(ptr_deref_804_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_804_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_804_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_817_addr_0
    process(ptr_deref_817_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_817_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_817_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_817_base_resize
    process(iNsTr_17_814) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_814;
      ov := iv(9 downto 0);
      ptr_deref_817_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_817_gather_scatter
    process(ptr_deref_817_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_817_data_0;
      ov(15 downto 0) := iv;
      iNsTr_18_818 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_817_root_address_inst
    process(ptr_deref_817_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_817_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_817_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_addr_0
    process(ptr_deref_880_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_880_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_base_resize
    process(scevgep_875) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep_875;
      ov := iv(9 downto 0);
      ptr_deref_880_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_gather_scatter
    process(iNsTr_30_878) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_30_878;
      ov(15 downto 0) := iv;
      ptr_deref_880_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_root_address_inst
    process(ptr_deref_880_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_880_root_address <= ov(9 downto 0);
      --
    end process;
    do_while_stmt_857_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_899_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_857_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_857_branch_req_0,
          ack0 => do_while_stmt_857_branch_ack_0,
          ack1 => do_while_stmt_857_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_776_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_775;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_776_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_776_branch_req_0,
          ack0 => if_stmt_776_branch_ack_0,
          ack1 => if_stmt_776_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_833_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_21_832;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_833_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_833_branch_req_0,
          ack0 => if_stmt_833_branch_ack_0,
          ack1 => if_stmt_833_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_900_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= bb_4_xx_x_crit_edgex_xloopexit_taken_896;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_900_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_900_branch_req_0,
          ack0 => if_stmt_900_branch_ack_0,
          ack1 => if_stmt_900_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u16_u16_843_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_12_792 & iNsTr_18_818;
      tmp_844 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_843_inst_req_0;
      ADD_u16_u16_843_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_843_inst_req_1;
      ADD_u16_u16_843_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u64_u64_768_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar7_744;
      indvarx_xnext8_769 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_768_inst_req_0;
      ADD_u64_u64_768_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_768_inst_req_1;
      ADD_u64_u64_768_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u64_u64_869_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar_859;
      tmp3_870 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_869_inst_req_0;
      ADD_u64_u64_869_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_869_inst_req_1;
      ADD_u64_u64_869_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u64_u64_887_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar_859;
      indvarx_xnext_888 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_887_inst_req_0;
      ADD_u64_u64_887_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_887_inst_req_1;
      ADD_u64_u64_887_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : EQ_u16_u1_831_inst 
    ApIntEq_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_12_792 & iNsTr_20_827;
      iNsTr_21_832 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_831_inst_req_0;
      EQ_u16_u1_831_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_831_inst_req_1;
      EQ_u16_u1_831_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_4_gI: SplitGuardInterface generic map(name => "ApIntEq_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : EQ_u64_u1_774_inst 
    ApIntEq_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnext8_769;
      exitcond_775 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_774_inst_req_0;
      EQ_u64_u1_774_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_774_inst_req_1;
      EQ_u64_u1_774_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_5_gI: SplitGuardInterface generic map(name => "ApIntEq_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : EQ_u64_u1_892_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnext_888 & tmp1_848;
      exitcond2_893 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_892_inst_req_0;
      EQ_u64_u1_892_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_892_inst_req_1;
      EQ_u64_u1_892_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- unary operator NOT_u1_u1_899_inst
    process(exitcond2_893) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", exitcond2_893, tmp_var);
      NOT_u1_u1_899_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (8) : SUB_u16_u16_826_inst 
    ApIntSub_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_824_wire_constant & iNsTr_18_818;
      iNsTr_20_827 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_826_inst_req_0;
      SUB_u16_u16_826_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_826_inst_req_1;
      SUB_u16_u16_826_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_8_gI: SplitGuardInterface generic map(name => "ApIntSub_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared load operator group (0) : ptr_deref_791_load_0 ptr_deref_804_load_0 ptr_deref_817_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_791_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_804_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_817_load_0_req_0;
      ptr_deref_791_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_804_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_817_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_791_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_804_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_817_load_0_req_1;
      ptr_deref_791_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_804_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_817_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_791_word_address_0 & ptr_deref_804_word_address_0 & ptr_deref_817_word_address_0;
      ptr_deref_791_data_0 <= data_out(47 downto 32);
      ptr_deref_804_data_0 <= data_out(31 downto 16);
      ptr_deref_817_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 10,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(9 downto 0),
          mtag => memory_space_8_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_ebbyNo_739_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ebbyNo_739_store_0_req_0;
      STORE_ebbyNo_739_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ebbyNo_739_store_0_req_1;
      STORE_ebbyNo_739_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ebbyNo_739_word_address_0;
      data_in <= STORE_ebbyNo_739_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_maxNitr_733_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_maxNitr_733_store_0_req_0;
      STORE_maxNitr_733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_maxNitr_733_store_0_req_1;
      STORE_maxNitr_733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_maxNitr_733_word_address_0;
      data_in <= STORE_maxNitr_733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_ncol_ind_819_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ncol_ind_819_store_0_req_0;
      STORE_ncol_ind_819_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ncol_ind_819_store_0_req_1;
      STORE_ncol_ind_819_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ncol_ind_819_word_address_0;
      data_in <= STORE_ncol_ind_819_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(0 downto 0),
          mdata => memory_space_10_sr_data(15 downto 0),
          mtag => memory_space_10_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : STORE_ncols_806_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_ncols_806_store_0_req_0;
      STORE_ncols_806_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_ncols_806_store_0_req_1;
      STORE_ncols_806_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ncols_806_word_address_0;
      data_in <= STORE_ncols_806_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(0 downto 0),
          mdata => memory_space_11_sr_data(15 downto 0),
          mtag => memory_space_11_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : STORE_nrows_793_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_nrows_793_store_0_req_0;
      STORE_nrows_793_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_nrows_793_store_0_req_1;
      STORE_nrows_793_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_nrows_793_word_address_0;
      data_in <= STORE_nrows_793_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_12_sr_req(0),
          mack => memory_space_12_sr_ack(0),
          maddr => memory_space_12_sr_addr(0 downto 0),
          mdata => memory_space_12_sr_data(15 downto 0),
          mtag => memory_space_12_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_12_sc_req(0),
          mack => memory_space_12_sc_ack(0),
          mtag => memory_space_12_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : STORE_rate_910_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_rate_910_store_0_req_0;
      STORE_rate_910_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_rate_910_store_0_req_1;
      STORE_rate_910_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_rate_910_word_address_0;
      data_in <= STORE_rate_910_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_13_sr_req(0),
          mack => memory_space_13_sr_ack(0),
          maddr => memory_space_13_sr_addr(0 downto 0),
          mdata => memory_space_13_sr_data(31 downto 0),
          mtag => memory_space_13_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_13_sc_req(0),
          mack => memory_space_13_sc_ack(0),
          mtag => memory_space_13_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_761_store_0 ptr_deref_880_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(19 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_761_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_880_store_0_req_0;
      ptr_deref_761_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_880_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_761_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_880_store_0_req_1;
      ptr_deref_761_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_880_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup6_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup6_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_761_word_address_0 & ptr_deref_880_word_address_0;
      data_in <= ptr_deref_761_data_0 & ptr_deref_880_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 10,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(9 downto 0),
          mdata => memory_space_8_sr_data(15 downto 0),
          mtag => memory_space_8_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_ebbyNo_in_737_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_ebbyNo_in_737_inst_req_0;
      RPIPE_ebbyNo_in_737_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_ebbyNo_in_737_inst_req_1;
      RPIPE_ebbyNo_in_737_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_4_738 <= data_out(31 downto 0);
      ebbyNo_in_read_0_gI: SplitGuardInterface generic map(name => "ebbyNo_in_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ebbyNo_in_read_0: InputPortRevised -- 
        generic map ( name => "ebbyNo_in_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ebbyNo_in_pipe_read_req(0),
          oack => ebbyNo_in_pipe_read_ack(0),
          odata => ebbyNo_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_matrix_in_758_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_matrix_in_758_inst_req_0;
      RPIPE_matrix_in_758_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_matrix_in_758_inst_req_1;
      RPIPE_matrix_in_758_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_8_759 <= data_out(15 downto 0);
      matrix_in_read_1_gI: SplitGuardInterface generic map(name => "matrix_in_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      matrix_in_read_1: InputPortRevised -- 
        generic map ( name => "matrix_in_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => matrix_in_pipe_read_req(1),
          oack => matrix_in_pipe_read_ack(1),
          odata => matrix_in_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_matrix_in_877_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_matrix_in_877_inst_req_0;
      RPIPE_matrix_in_877_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_matrix_in_877_inst_req_1;
      RPIPE_matrix_in_877_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_30_878 <= data_out(15 downto 0);
      matrix_in_read_2_gI: SplitGuardInterface generic map(name => "matrix_in_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      matrix_in_read_2: InputPortRevised -- 
        generic map ( name => "matrix_in_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => matrix_in_pipe_read_req(0),
          oack => matrix_in_pipe_read_ack(0),
          odata => matrix_in_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_maxNitr_in_731_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_maxNitr_in_731_inst_req_0;
      RPIPE_maxNitr_in_731_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_maxNitr_in_731_inst_req_1;
      RPIPE_maxNitr_in_731_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_1_732 <= data_out(15 downto 0);
      maxNitr_in_read_3_gI: SplitGuardInterface generic map(name => "maxNitr_in_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxNitr_in_read_3: InputPortRevised -- 
        generic map ( name => "maxNitr_in_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxNitr_in_pipe_read_req(0),
          oack => maxNitr_in_pipe_read_ack(0),
          odata => maxNitr_in_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_rate_in_908_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_rate_in_908_inst_req_0;
      RPIPE_rate_in_908_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_rate_in_908_inst_req_1;
      RPIPE_rate_in_908_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_24_909 <= data_out(31 downto 0);
      rate_in_read_4_gI: SplitGuardInterface generic map(name => "rate_in_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      rate_in_read_4: InputPortRevised -- 
        generic map ( name => "rate_in_read_4", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => rate_in_pipe_read_req(0),
          oack => rate_in_pipe_read_ack(0),
          odata => rate_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- 
  end Block; -- data_path
  -- 
end initInputs_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity minSumDecode is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_11_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_11_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_11_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_11_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_11_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_11_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(9 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_10_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_12_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_12_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_12_lr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_12_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_12_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_12_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_12_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_13_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_13_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_13_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_13_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_13_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_13_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_13_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_9_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_9_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(5 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
    code_block_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    code_block_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    code_block_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    code_block_decoded_pipe_write_req : out  std_logic_vector(0 downto 0);
    code_block_decoded_pipe_write_ack : in   std_logic_vector(0 downto 0);
    code_block_decoded_pipe_write_data : out  std_logic_vector(31 downto 0);
    nitr_required_pipe_write_req : out  std_logic_vector(0 downto 0);
    nitr_required_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nitr_required_pipe_write_data : out  std_logic_vector(15 downto 0);
    checkNodeComputeEngine_call_reqs : out  std_logic_vector(0 downto 0);
    checkNodeComputeEngine_call_acks : in   std_logic_vector(0 downto 0);
    checkNodeComputeEngine_call_tag  :  out  std_logic_vector(0 downto 0);
    checkNodeComputeEngine_return_reqs : out  std_logic_vector(0 downto 0);
    checkNodeComputeEngine_return_acks : in   std_logic_vector(0 downto 0);
    checkNodeComputeEngine_return_tag :  in   std_logic_vector(0 downto 0);
    initInputs_call_reqs : out  std_logic_vector(0 downto 0);
    initInputs_call_acks : in   std_logic_vector(0 downto 0);
    initInputs_call_tag  :  out  std_logic_vector(0 downto 0);
    initInputs_return_reqs : out  std_logic_vector(0 downto 0);
    initInputs_return_acks : in   std_logic_vector(0 downto 0);
    initInputs_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity minSumDecode;
architecture minSumDecode_arch of minSumDecode is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal minSumDecode_CP_6680_start: Boolean;
  signal minSumDecode_CP_6680_symbol: Boolean;
  -- volatile/operator module components. 
  component checkNodeComputeEngine is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_9_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_9_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_9_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_9_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_12_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_12_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_12_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component initInputs is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_11_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_12_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_12_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_12_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_12_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_13_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_13_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_13_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_13_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sc_tag :  in  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      matrix_in_pipe_read_req : out  std_logic_vector(1 downto 0);
      matrix_in_pipe_read_ack : in   std_logic_vector(1 downto 0);
      matrix_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal addr_of_1520_final_reg_req_0 : boolean;
  signal addr_of_1520_final_reg_ack_0 : boolean;
  signal addr_of_1520_final_reg_req_1 : boolean;
  signal addr_of_1520_final_reg_ack_1 : boolean;
  signal call_stmt_1356_call_req_0 : boolean;
  signal call_stmt_1356_call_ack_0 : boolean;
  signal call_stmt_1356_call_req_1 : boolean;
  signal call_stmt_1356_call_ack_1 : boolean;
  signal LOAD_ncols_1358_load_0_req_0 : boolean;
  signal LOAD_ncols_1358_load_0_ack_0 : boolean;
  signal LOAD_ncols_1358_load_0_req_1 : boolean;
  signal LOAD_ncols_1358_load_0_ack_1 : boolean;
  signal EQ_u16_u1_1364_inst_req_0 : boolean;
  signal EQ_u16_u1_1364_inst_ack_0 : boolean;
  signal EQ_u16_u1_1364_inst_req_1 : boolean;
  signal EQ_u16_u1_1364_inst_ack_1 : boolean;
  signal if_stmt_1366_branch_req_0 : boolean;
  signal if_stmt_1366_branch_ack_1 : boolean;
  signal if_stmt_1366_branch_ack_0 : boolean;
  signal do_while_stmt_1381_branch_req_0 : boolean;
  signal phi_stmt_1383_req_0 : boolean;
  signal phi_stmt_1383_req_1 : boolean;
  signal phi_stmt_1383_ack_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal iNsTr_13_at_entry_1375_1387_buf_req_0 : boolean;
  signal iNsTr_13_at_entry_1375_1387_buf_ack_0 : boolean;
  signal iNsTr_13_at_entry_1375_1387_buf_req_1 : boolean;
  signal iNsTr_13_at_entry_1375_1387_buf_ack_1 : boolean;
  signal ptr_deref_1805_load_0_req_1 : boolean;
  signal ADD_u8_u8_1393_inst_req_0 : boolean;
  signal ADD_u8_u8_1393_inst_ack_0 : boolean;
  signal ADD_u8_u8_1393_inst_req_1 : boolean;
  signal ADD_u8_u8_1393_inst_ack_1 : boolean;
  signal ADD_u8_u8_1399_inst_req_0 : boolean;
  signal ADD_u8_u8_1399_inst_ack_0 : boolean;
  signal ADD_u8_u8_1399_inst_req_1 : boolean;
  signal ADD_u8_u8_1399_inst_ack_1 : boolean;
  signal RPIPE_code_block_in_1402_inst_req_0 : boolean;
  signal RPIPE_code_block_in_1402_inst_ack_0 : boolean;
  signal RPIPE_code_block_in_1402_inst_req_1 : boolean;
  signal RPIPE_code_block_in_1402_inst_ack_1 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal addr_of_1801_final_reg_req_1 : boolean;
  signal ptr_deref_1805_load_0_ack_1 : boolean;
  signal addr_of_1411_final_reg_req_0 : boolean;
  signal addr_of_1411_final_reg_ack_0 : boolean;
  signal addr_of_1411_final_reg_req_1 : boolean;
  signal addr_of_1411_final_reg_ack_1 : boolean;
  signal addr_of_1801_final_reg_ack_1 : boolean;
  signal ptr_deref_1414_store_0_req_0 : boolean;
  signal ptr_deref_1414_store_0_ack_0 : boolean;
  signal ptr_deref_1414_store_0_req_1 : boolean;
  signal ptr_deref_1414_store_0_ack_1 : boolean;
  signal addr_of_1801_final_reg_ack_0 : boolean;
  signal type_cast_1419_inst_req_0 : boolean;
  signal type_cast_1419_inst_ack_0 : boolean;
  signal ptr_deref_1805_load_0_req_0 : boolean;
  signal type_cast_1419_inst_req_1 : boolean;
  signal type_cast_1419_inst_ack_1 : boolean;
  signal ptr_deref_1805_load_0_ack_0 : boolean;
  signal addr_of_1801_final_reg_req_0 : boolean;
  signal LOAD_ncols_1422_load_0_req_0 : boolean;
  signal LOAD_ncols_1422_load_0_ack_0 : boolean;
  signal LOAD_ncols_1422_load_0_req_1 : boolean;
  signal LOAD_ncols_1422_load_0_ack_1 : boolean;
  signal type_cast_1426_inst_req_0 : boolean;
  signal type_cast_1426_inst_ack_0 : boolean;
  signal type_cast_1426_inst_req_1 : boolean;
  signal type_cast_1426_inst_ack_1 : boolean;
  signal ULT_u32_u1_1431_inst_req_0 : boolean;
  signal ULT_u32_u1_1431_inst_ack_0 : boolean;
  signal ULT_u32_u1_1431_inst_req_1 : boolean;
  signal ULT_u32_u1_1431_inst_ack_1 : boolean;
  signal NOT_u1_u1_1435_inst_req_0 : boolean;
  signal NOT_u1_u1_1435_inst_ack_0 : boolean;
  signal NOT_u1_u1_1435_inst_req_1 : boolean;
  signal NOT_u1_u1_1435_inst_ack_1 : boolean;
  signal do_while_stmt_1381_branch_ack_0 : boolean;
  signal do_while_stmt_1381_branch_ack_1 : boolean;
  signal if_stmt_1439_branch_req_0 : boolean;
  signal if_stmt_1439_branch_ack_1 : boolean;
  signal if_stmt_1439_branch_ack_0 : boolean;
  signal EQ_u16_u1_1453_inst_req_0 : boolean;
  signal EQ_u16_u1_1453_inst_ack_0 : boolean;
  signal EQ_u16_u1_1453_inst_req_1 : boolean;
  signal EQ_u16_u1_1453_inst_ack_1 : boolean;
  signal if_stmt_1455_branch_req_0 : boolean;
  signal if_stmt_1455_branch_ack_1 : boolean;
  signal if_stmt_1455_branch_ack_0 : boolean;
  signal LOAD_ebbyNo_1463_load_0_req_0 : boolean;
  signal LOAD_ebbyNo_1463_load_0_ack_0 : boolean;
  signal LOAD_ebbyNo_1463_load_0_req_1 : boolean;
  signal LOAD_ebbyNo_1463_load_0_ack_1 : boolean;
  signal LOAD_rate_1466_load_0_req_0 : boolean;
  signal LOAD_rate_1466_load_0_ack_0 : boolean;
  signal LOAD_rate_1466_load_0_req_1 : boolean;
  signal LOAD_rate_1466_load_0_ack_1 : boolean;
  signal MUL_f32_f32_1471_inst_req_0 : boolean;
  signal MUL_f32_f32_1471_inst_ack_0 : boolean;
  signal MUL_f32_f32_1471_inst_req_1 : boolean;
  signal MUL_f32_f32_1471_inst_ack_1 : boolean;
  signal UGT_u16_u1_1477_inst_req_0 : boolean;
  signal UGT_u16_u1_1477_inst_ack_0 : boolean;
  signal UGT_u16_u1_1477_inst_req_1 : boolean;
  signal UGT_u16_u1_1477_inst_ack_1 : boolean;
  signal ADD_u16_u16_1483_inst_req_0 : boolean;
  signal ADD_u16_u16_1483_inst_ack_0 : boolean;
  signal ADD_u16_u16_1483_inst_req_1 : boolean;
  signal ADD_u16_u16_1483_inst_ack_1 : boolean;
  signal type_cast_1487_inst_req_0 : boolean;
  signal type_cast_1487_inst_ack_0 : boolean;
  signal type_cast_1487_inst_req_1 : boolean;
  signal type_cast_1487_inst_ack_1 : boolean;
  signal ADD_u64_u64_1493_inst_req_0 : boolean;
  signal ADD_u64_u64_1493_inst_ack_0 : boolean;
  signal ADD_u64_u64_1493_inst_req_1 : boolean;
  signal ADD_u64_u64_1493_inst_ack_1 : boolean;
  signal MUX_1500_inst_req_0 : boolean;
  signal MUX_1500_inst_ack_0 : boolean;
  signal MUX_1500_inst_req_1 : boolean;
  signal MUX_1500_inst_ack_1 : boolean;
  signal addr_of_1515_final_reg_req_0 : boolean;
  signal addr_of_1515_final_reg_ack_0 : boolean;
  signal addr_of_1515_final_reg_req_1 : boolean;
  signal addr_of_1515_final_reg_ack_1 : boolean;
  signal ptr_deref_1524_load_0_req_0 : boolean;
  signal ptr_deref_1524_load_0_ack_0 : boolean;
  signal ptr_deref_1524_load_0_req_1 : boolean;
  signal ptr_deref_1524_load_0_ack_1 : boolean;
  signal MUL_f32_f32_1530_inst_req_0 : boolean;
  signal MUL_f32_f32_1530_inst_ack_0 : boolean;
  signal MUL_f32_f32_1530_inst_req_1 : boolean;
  signal MUL_f32_f32_1530_inst_ack_1 : boolean;
  signal MUL_f32_f32_1535_inst_req_0 : boolean;
  signal MUL_f32_f32_1535_inst_ack_0 : boolean;
  signal MUL_f32_f32_1535_inst_req_1 : boolean;
  signal MUL_f32_f32_1535_inst_ack_1 : boolean;
  signal ptr_deref_1538_store_0_req_0 : boolean;
  signal ptr_deref_1538_store_0_ack_0 : boolean;
  signal ptr_deref_1538_store_0_req_1 : boolean;
  signal ptr_deref_1538_store_0_ack_1 : boolean;
  signal ADD_u64_u64_1545_inst_req_0 : boolean;
  signal ADD_u64_u64_1545_inst_ack_0 : boolean;
  signal ADD_u64_u64_1545_inst_req_1 : boolean;
  signal ADD_u64_u64_1545_inst_ack_1 : boolean;
  signal EQ_u64_u1_1550_inst_req_0 : boolean;
  signal EQ_u64_u1_1550_inst_ack_0 : boolean;
  signal EQ_u64_u1_1550_inst_req_1 : boolean;
  signal EQ_u64_u1_1550_inst_ack_1 : boolean;
  signal if_stmt_1552_branch_req_0 : boolean;
  signal if_stmt_1552_branch_ack_1 : boolean;
  signal if_stmt_1552_branch_ack_0 : boolean;
  signal LOAD_ncol_ind_1573_load_0_req_0 : boolean;
  signal LOAD_ncol_ind_1573_load_0_ack_0 : boolean;
  signal LOAD_ncol_ind_1573_load_0_req_1 : boolean;
  signal LOAD_ncol_ind_1573_load_0_ack_1 : boolean;
  signal EQ_u16_u1_1579_inst_req_0 : boolean;
  signal EQ_u16_u1_1579_inst_ack_0 : boolean;
  signal EQ_u16_u1_1579_inst_req_1 : boolean;
  signal EQ_u16_u1_1579_inst_ack_1 : boolean;
  signal if_stmt_1581_branch_req_0 : boolean;
  signal if_stmt_1581_branch_ack_1 : boolean;
  signal if_stmt_1581_branch_ack_0 : boolean;
  signal UGT_u16_u1_1592_inst_req_0 : boolean;
  signal UGT_u16_u1_1592_inst_ack_0 : boolean;
  signal UGT_u16_u1_1592_inst_req_1 : boolean;
  signal UGT_u16_u1_1592_inst_ack_1 : boolean;
  signal ADD_u16_u16_1598_inst_req_0 : boolean;
  signal ADD_u16_u16_1598_inst_ack_0 : boolean;
  signal ADD_u16_u16_1598_inst_req_1 : boolean;
  signal ADD_u16_u16_1598_inst_ack_1 : boolean;
  signal type_cast_1602_inst_req_0 : boolean;
  signal type_cast_1602_inst_ack_0 : boolean;
  signal type_cast_1602_inst_req_1 : boolean;
  signal type_cast_1602_inst_ack_1 : boolean;
  signal ADD_u64_u64_1608_inst_req_0 : boolean;
  signal ADD_u64_u64_1608_inst_ack_0 : boolean;
  signal ADD_u64_u64_1608_inst_req_1 : boolean;
  signal ADD_u64_u64_1608_inst_ack_1 : boolean;
  signal MUX_1615_inst_req_0 : boolean;
  signal MUX_1615_inst_ack_0 : boolean;
  signal MUX_1615_inst_req_1 : boolean;
  signal MUX_1615_inst_ack_1 : boolean;
  signal addr_of_1630_final_reg_req_0 : boolean;
  signal addr_of_1630_final_reg_ack_0 : boolean;
  signal addr_of_1630_final_reg_req_1 : boolean;
  signal addr_of_1630_final_reg_ack_1 : boolean;
  signal ADD_u64_u64_1636_inst_req_0 : boolean;
  signal ADD_u64_u64_1636_inst_ack_0 : boolean;
  signal ADD_u64_u64_1636_inst_req_1 : boolean;
  signal ADD_u64_u64_1636_inst_ack_1 : boolean;
  signal addr_of_1641_final_reg_req_0 : boolean;
  signal addr_of_1641_final_reg_ack_0 : boolean;
  signal addr_of_1641_final_reg_req_1 : boolean;
  signal addr_of_1641_final_reg_ack_1 : boolean;
  signal ptr_deref_1645_load_0_req_0 : boolean;
  signal ptr_deref_1645_load_0_ack_0 : boolean;
  signal ptr_deref_1645_load_0_req_1 : boolean;
  signal ptr_deref_1645_load_0_ack_1 : boolean;
  signal ADD_u16_u16_1651_inst_req_0 : boolean;
  signal ADD_u16_u16_1651_inst_ack_0 : boolean;
  signal ADD_u16_u16_1651_inst_req_1 : boolean;
  signal ADD_u16_u16_1651_inst_ack_1 : boolean;
  signal type_cast_1655_inst_req_0 : boolean;
  signal type_cast_1655_inst_ack_0 : boolean;
  signal type_cast_1655_inst_req_1 : boolean;
  signal type_cast_1655_inst_ack_1 : boolean;
  signal EQ_u64_u1_2030_inst_ack_1 : boolean;
  signal addr_of_1660_final_reg_req_0 : boolean;
  signal addr_of_1660_final_reg_ack_0 : boolean;
  signal addr_of_1660_final_reg_req_1 : boolean;
  signal addr_of_1660_final_reg_ack_1 : boolean;
  signal ptr_deref_1664_load_0_req_0 : boolean;
  signal ptr_deref_1664_load_0_ack_0 : boolean;
  signal ptr_deref_1664_load_0_req_1 : boolean;
  signal ptr_deref_1664_load_0_ack_1 : boolean;
  signal EQ_u64_u1_2030_inst_ack_0 : boolean;
  signal if_stmt_2054_branch_req_0 : boolean;
  signal ptr_deref_1667_store_0_req_0 : boolean;
  signal ptr_deref_1667_store_0_ack_0 : boolean;
  signal ptr_deref_1667_store_0_req_1 : boolean;
  signal ptr_deref_1667_store_0_ack_1 : boolean;
  signal ADD_u64_u64_1674_inst_req_0 : boolean;
  signal ADD_u64_u64_1674_inst_ack_0 : boolean;
  signal ADD_u64_u64_1674_inst_req_1 : boolean;
  signal ADD_u64_u64_1674_inst_ack_1 : boolean;
  signal EQ_u64_u1_1679_inst_req_0 : boolean;
  signal EQ_u64_u1_1679_inst_ack_0 : boolean;
  signal EQ_u64_u1_1679_inst_req_1 : boolean;
  signal EQ_u64_u1_1679_inst_ack_1 : boolean;
  signal if_stmt_2054_branch_ack_1 : boolean;
  signal if_stmt_1681_branch_req_0 : boolean;
  signal EQ_u64_u1_2030_inst_req_1 : boolean;
  signal if_stmt_1681_branch_ack_1 : boolean;
  signal if_stmt_1681_branch_ack_0 : boolean;
  signal ADD_u16_u16_1724_inst_req_0 : boolean;
  signal ADD_u16_u16_1724_inst_ack_0 : boolean;
  signal LOAD_ncols_2046_load_0_req_0 : boolean;
  signal ADD_u16_u16_1724_inst_req_1 : boolean;
  signal ADD_u16_u16_1724_inst_ack_1 : boolean;
  signal LOAD_maxNitr_1727_load_0_req_0 : boolean;
  signal LOAD_maxNitr_1727_load_0_ack_0 : boolean;
  signal LOAD_ncols_2046_load_0_ack_0 : boolean;
  signal LOAD_maxNitr_1727_load_0_req_1 : boolean;
  signal LOAD_maxNitr_1727_load_0_ack_1 : boolean;
  signal ULT_u16_u1_1732_inst_req_0 : boolean;
  signal ULT_u16_u1_1732_inst_ack_0 : boolean;
  signal ULT_u16_u1_1732_inst_req_1 : boolean;
  signal ULT_u16_u1_1732_inst_ack_1 : boolean;
  signal if_stmt_1734_branch_req_0 : boolean;
  signal if_stmt_1734_branch_ack_1 : boolean;
  signal if_stmt_1734_branch_ack_0 : boolean;
  signal EQ_u64_u1_2030_inst_req_0 : boolean;
  signal EQ_u16_u1_1745_inst_req_0 : boolean;
  signal EQ_u16_u1_1745_inst_ack_0 : boolean;
  signal EQ_u16_u1_1745_inst_req_1 : boolean;
  signal EQ_u16_u1_1745_inst_ack_1 : boolean;
  signal if_stmt_1747_branch_req_0 : boolean;
  signal if_stmt_1747_branch_ack_1 : boolean;
  signal if_stmt_1747_branch_ack_0 : boolean;
  signal UGT_u16_u1_1758_inst_req_0 : boolean;
  signal UGT_u16_u1_1758_inst_ack_0 : boolean;
  signal UGT_u16_u1_1758_inst_req_1 : boolean;
  signal UGT_u16_u1_1758_inst_ack_1 : boolean;
  signal ADD_u16_u16_1764_inst_req_0 : boolean;
  signal ADD_u16_u16_1764_inst_ack_0 : boolean;
  signal ADD_u16_u16_1764_inst_req_1 : boolean;
  signal ADD_u16_u16_1764_inst_ack_1 : boolean;
  signal type_cast_1768_inst_req_0 : boolean;
  signal type_cast_1768_inst_ack_0 : boolean;
  signal type_cast_1768_inst_req_1 : boolean;
  signal type_cast_1768_inst_ack_1 : boolean;
  signal ADD_u64_u64_1774_inst_req_0 : boolean;
  signal ADD_u64_u64_1774_inst_ack_0 : boolean;
  signal ADD_u64_u64_1774_inst_req_1 : boolean;
  signal ADD_u64_u64_1774_inst_ack_1 : boolean;
  signal MUX_1781_inst_req_0 : boolean;
  signal MUX_1781_inst_ack_0 : boolean;
  signal MUX_1781_inst_req_1 : boolean;
  signal MUX_1781_inst_ack_1 : boolean;
  signal addr_of_1796_final_reg_req_0 : boolean;
  signal addr_of_1796_final_reg_ack_0 : boolean;
  signal addr_of_1796_final_reg_req_1 : boolean;
  signal addr_of_1796_final_reg_ack_1 : boolean;
  signal ptr_deref_1808_store_0_req_0 : boolean;
  signal ptr_deref_1808_store_0_ack_0 : boolean;
  signal ptr_deref_1808_store_0_req_1 : boolean;
  signal ptr_deref_1808_store_0_ack_1 : boolean;
  signal ADD_u64_u64_1815_inst_req_0 : boolean;
  signal ADD_u64_u64_1815_inst_ack_0 : boolean;
  signal ADD_u64_u64_1815_inst_req_1 : boolean;
  signal ADD_u64_u64_1815_inst_ack_1 : boolean;
  signal EQ_u64_u1_1820_inst_req_0 : boolean;
  signal EQ_u64_u1_1820_inst_ack_0 : boolean;
  signal EQ_u64_u1_1820_inst_req_1 : boolean;
  signal EQ_u64_u1_1820_inst_ack_1 : boolean;
  signal if_stmt_1822_branch_req_0 : boolean;
  signal if_stmt_1822_branch_ack_1 : boolean;
  signal if_stmt_1822_branch_ack_0 : boolean;
  signal EQ_u16_u1_1835_inst_req_0 : boolean;
  signal EQ_u16_u1_1835_inst_ack_0 : boolean;
  signal EQ_u16_u1_1835_inst_req_1 : boolean;
  signal EQ_u16_u1_1835_inst_ack_1 : boolean;
  signal if_stmt_1837_branch_req_0 : boolean;
  signal if_stmt_1837_branch_ack_1 : boolean;
  signal if_stmt_1837_branch_ack_0 : boolean;
  signal UGT_u16_u1_1848_inst_req_0 : boolean;
  signal UGT_u16_u1_1848_inst_ack_0 : boolean;
  signal UGT_u16_u1_1848_inst_req_1 : boolean;
  signal UGT_u16_u1_1848_inst_ack_1 : boolean;
  signal ADD_u16_u16_1854_inst_req_0 : boolean;
  signal ADD_u16_u16_1854_inst_ack_0 : boolean;
  signal ADD_u16_u16_1854_inst_req_1 : boolean;
  signal ADD_u16_u16_1854_inst_ack_1 : boolean;
  signal type_cast_1858_inst_req_0 : boolean;
  signal type_cast_1858_inst_ack_0 : boolean;
  signal type_cast_1858_inst_req_1 : boolean;
  signal type_cast_1858_inst_ack_1 : boolean;
  signal ADD_u64_u64_1864_inst_req_0 : boolean;
  signal ADD_u64_u64_1864_inst_ack_0 : boolean;
  signal ADD_u64_u64_1864_inst_req_1 : boolean;
  signal ADD_u64_u64_1864_inst_ack_1 : boolean;
  signal MUX_1871_inst_req_0 : boolean;
  signal MUX_1871_inst_ack_0 : boolean;
  signal MUX_1871_inst_req_1 : boolean;
  signal MUX_1871_inst_ack_1 : boolean;
  signal addr_of_1886_final_reg_req_0 : boolean;
  signal addr_of_1886_final_reg_ack_0 : boolean;
  signal addr_of_1886_final_reg_req_1 : boolean;
  signal addr_of_1886_final_reg_ack_1 : boolean;
  signal ptr_deref_1889_store_0_req_0 : boolean;
  signal ptr_deref_1889_store_0_ack_0 : boolean;
  signal ptr_deref_1889_store_0_req_1 : boolean;
  signal ptr_deref_1889_store_0_ack_1 : boolean;
  signal ADD_u64_u64_1897_inst_req_0 : boolean;
  signal ADD_u64_u64_1897_inst_ack_0 : boolean;
  signal ADD_u64_u64_1897_inst_req_1 : boolean;
  signal ADD_u64_u64_1897_inst_ack_1 : boolean;
  signal EQ_u64_u1_1902_inst_req_0 : boolean;
  signal EQ_u64_u1_1902_inst_ack_0 : boolean;
  signal EQ_u64_u1_1902_inst_req_1 : boolean;
  signal EQ_u64_u1_1902_inst_ack_1 : boolean;
  signal if_stmt_1904_branch_req_0 : boolean;
  signal if_stmt_1904_branch_ack_1 : boolean;
  signal if_stmt_1904_branch_ack_0 : boolean;
  signal call_stmt_1913_call_req_0 : boolean;
  signal call_stmt_1913_call_ack_0 : boolean;
  signal call_stmt_1913_call_req_1 : boolean;
  signal call_stmt_1913_call_ack_1 : boolean;
  signal LOAD_ncol_ind_1915_load_0_req_0 : boolean;
  signal LOAD_ncol_ind_1915_load_0_ack_0 : boolean;
  signal LOAD_ncol_ind_1915_load_0_req_1 : boolean;
  signal LOAD_ncol_ind_1915_load_0_ack_1 : boolean;
  signal EQ_u16_u1_1921_inst_req_0 : boolean;
  signal EQ_u16_u1_1921_inst_ack_0 : boolean;
  signal EQ_u16_u1_1921_inst_req_1 : boolean;
  signal EQ_u16_u1_1921_inst_ack_1 : boolean;
  signal if_stmt_1923_branch_req_0 : boolean;
  signal if_stmt_1923_branch_ack_1 : boolean;
  signal if_stmt_1923_branch_ack_0 : boolean;
  signal UGT_u16_u1_1934_inst_req_0 : boolean;
  signal UGT_u16_u1_1934_inst_ack_0 : boolean;
  signal UGT_u16_u1_1934_inst_req_1 : boolean;
  signal UGT_u16_u1_1934_inst_ack_1 : boolean;
  signal ADD_u16_u16_1940_inst_req_0 : boolean;
  signal ADD_u16_u16_1940_inst_ack_0 : boolean;
  signal ADD_u16_u16_1940_inst_req_1 : boolean;
  signal ADD_u16_u16_1940_inst_ack_1 : boolean;
  signal type_cast_1944_inst_req_0 : boolean;
  signal type_cast_1944_inst_ack_0 : boolean;
  signal type_cast_1944_inst_req_1 : boolean;
  signal type_cast_1944_inst_ack_1 : boolean;
  signal ADD_u64_u64_1950_inst_req_0 : boolean;
  signal ADD_u64_u64_1950_inst_ack_0 : boolean;
  signal ADD_u64_u64_1950_inst_req_1 : boolean;
  signal ADD_u64_u64_1950_inst_ack_1 : boolean;
  signal MUX_1957_inst_req_0 : boolean;
  signal MUX_1957_inst_ack_0 : boolean;
  signal MUX_1957_inst_req_1 : boolean;
  signal MUX_1957_inst_ack_1 : boolean;
  signal STORE_is_decoded_2041_store_0_ack_1 : boolean;
  signal addr_of_1972_final_reg_req_0 : boolean;
  signal addr_of_1972_final_reg_ack_0 : boolean;
  signal STORE_is_decoded_2041_store_0_req_1 : boolean;
  signal addr_of_1972_final_reg_req_1 : boolean;
  signal addr_of_1972_final_reg_ack_1 : boolean;
  signal ADD_u64_u64_1978_inst_req_0 : boolean;
  signal ADD_u64_u64_1978_inst_ack_0 : boolean;
  signal ADD_u64_u64_1978_inst_req_1 : boolean;
  signal ADD_u64_u64_1978_inst_ack_1 : boolean;
  signal if_stmt_2032_branch_req_0 : boolean;
  signal if_stmt_2054_branch_ack_0 : boolean;
  signal STORE_is_decoded_2041_store_0_ack_0 : boolean;
  signal addr_of_1983_final_reg_req_0 : boolean;
  signal addr_of_1983_final_reg_ack_0 : boolean;
  signal STORE_is_decoded_2041_store_0_req_0 : boolean;
  signal addr_of_1983_final_reg_req_1 : boolean;
  signal addr_of_1983_final_reg_ack_1 : boolean;
  signal EQ_u16_u1_2052_inst_ack_1 : boolean;
  signal EQ_u16_u1_2052_inst_req_1 : boolean;
  signal ptr_deref_1987_load_0_req_0 : boolean;
  signal ptr_deref_1987_load_0_ack_0 : boolean;
  signal ptr_deref_1987_load_0_req_1 : boolean;
  signal ptr_deref_1987_load_0_ack_1 : boolean;
  signal EQ_u16_u1_2052_inst_ack_0 : boolean;
  signal EQ_u16_u1_2052_inst_req_0 : boolean;
  signal ADD_u16_u16_1993_inst_req_0 : boolean;
  signal ADD_u16_u16_1993_inst_ack_0 : boolean;
  signal ADD_u16_u16_1993_inst_req_1 : boolean;
  signal ADD_u16_u16_1993_inst_ack_1 : boolean;
  signal ptr_deref_1997_load_0_req_0 : boolean;
  signal ptr_deref_1997_load_0_ack_0 : boolean;
  signal if_stmt_2032_branch_ack_0 : boolean;
  signal ptr_deref_1997_load_0_req_1 : boolean;
  signal ptr_deref_1997_load_0_ack_1 : boolean;
  signal if_stmt_2032_branch_ack_1 : boolean;
  signal LOAD_ncols_2046_load_0_ack_1 : boolean;
  signal type_cast_2001_inst_req_0 : boolean;
  signal type_cast_2001_inst_ack_0 : boolean;
  signal type_cast_2001_inst_req_1 : boolean;
  signal type_cast_2001_inst_ack_1 : boolean;
  signal LOAD_ncols_2046_load_0_req_1 : boolean;
  signal ADD_u64_u64_2394_inst_ack_1 : boolean;
  signal ADD_u64_u64_2380_inst_ack_1 : boolean;
  signal addr_of_2006_final_reg_req_0 : boolean;
  signal addr_of_2006_final_reg_ack_0 : boolean;
  signal addr_of_2006_final_reg_req_1 : boolean;
  signal addr_of_2006_final_reg_ack_1 : boolean;
  signal type_cast_2389_inst_req_0 : boolean;
  signal type_cast_2389_inst_ack_0 : boolean;
  signal ADD_u64_u64_2380_inst_ack_0 : boolean;
  signal ptr_deref_2010_load_0_req_0 : boolean;
  signal ptr_deref_2010_load_0_ack_0 : boolean;
  signal ADD_u64_u64_2380_inst_req_0 : boolean;
  signal ptr_deref_2010_load_0_req_1 : boolean;
  signal ptr_deref_2010_load_0_ack_1 : boolean;
  signal ADD_u64_u64_2394_inst_req_1 : boolean;
  signal ADD_f32_f32_2015_inst_req_0 : boolean;
  signal ADD_f32_f32_2015_inst_ack_0 : boolean;
  signal ADD_f32_f32_2015_inst_req_1 : boolean;
  signal ADD_f32_f32_2015_inst_ack_1 : boolean;
  signal ptr_deref_2018_store_0_req_0 : boolean;
  signal ptr_deref_2018_store_0_ack_0 : boolean;
  signal ptr_deref_2018_store_0_req_1 : boolean;
  signal ptr_deref_2018_store_0_ack_1 : boolean;
  signal ADD_u64_u64_2025_inst_req_0 : boolean;
  signal ADD_u64_u64_2025_inst_ack_0 : boolean;
  signal ADD_u64_u64_2025_inst_req_1 : boolean;
  signal ADD_u64_u64_2025_inst_ack_1 : boolean;
  signal STORE_Nitr_required_2066_store_0_req_0 : boolean;
  signal STORE_Nitr_required_2066_store_0_ack_0 : boolean;
  signal STORE_Nitr_required_2066_store_0_req_1 : boolean;
  signal STORE_Nitr_required_2066_store_0_ack_1 : boolean;
  signal UGT_u16_u1_2075_inst_req_0 : boolean;
  signal UGT_u16_u1_2075_inst_ack_0 : boolean;
  signal UGT_u16_u1_2075_inst_req_1 : boolean;
  signal UGT_u16_u1_2075_inst_ack_1 : boolean;
  signal ADD_u16_u16_2081_inst_req_0 : boolean;
  signal ADD_u16_u16_2081_inst_ack_0 : boolean;
  signal ADD_u16_u16_2081_inst_req_1 : boolean;
  signal ADD_u16_u16_2081_inst_ack_1 : boolean;
  signal type_cast_2085_inst_req_0 : boolean;
  signal type_cast_2085_inst_ack_0 : boolean;
  signal type_cast_2085_inst_req_1 : boolean;
  signal type_cast_2085_inst_ack_1 : boolean;
  signal ADD_u64_u64_2091_inst_req_0 : boolean;
  signal ADD_u64_u64_2091_inst_ack_0 : boolean;
  signal ADD_u64_u64_2091_inst_req_1 : boolean;
  signal ADD_u64_u64_2091_inst_ack_1 : boolean;
  signal MUX_2098_inst_req_0 : boolean;
  signal MUX_2098_inst_ack_0 : boolean;
  signal MUX_2098_inst_req_1 : boolean;
  signal MUX_2098_inst_ack_1 : boolean;
  signal addr_of_2120_final_reg_req_0 : boolean;
  signal addr_of_2120_final_reg_ack_0 : boolean;
  signal addr_of_2120_final_reg_req_1 : boolean;
  signal addr_of_2120_final_reg_ack_1 : boolean;
  signal addr_of_2125_final_reg_req_0 : boolean;
  signal addr_of_2125_final_reg_ack_0 : boolean;
  signal addr_of_2125_final_reg_req_1 : boolean;
  signal addr_of_2125_final_reg_ack_1 : boolean;
  signal ptr_deref_2129_load_0_req_0 : boolean;
  signal ptr_deref_2129_load_0_ack_0 : boolean;
  signal ptr_deref_2129_load_0_req_1 : boolean;
  signal ptr_deref_2129_load_0_ack_1 : boolean;
  signal type_cast_2133_inst_req_0 : boolean;
  signal type_cast_2133_inst_ack_0 : boolean;
  signal type_cast_2133_inst_req_1 : boolean;
  signal type_cast_2133_inst_ack_1 : boolean;
  signal SGT_f64_u1_2139_inst_req_0 : boolean;
  signal SGT_f64_u1_2139_inst_ack_0 : boolean;
  signal SGT_f64_u1_2139_inst_req_1 : boolean;
  signal SGT_f64_u1_2139_inst_ack_1 : boolean;
  signal if_stmt_2141_branch_req_0 : boolean;
  signal if_stmt_2141_branch_ack_1 : boolean;
  signal if_stmt_2141_branch_ack_0 : boolean;
  signal ptr_deref_2150_load_0_req_0 : boolean;
  signal ptr_deref_2150_load_0_ack_0 : boolean;
  signal ptr_deref_2150_load_0_req_1 : boolean;
  signal ptr_deref_2150_load_0_ack_1 : boolean;
  signal type_cast_2154_inst_req_0 : boolean;
  signal type_cast_2154_inst_ack_0 : boolean;
  signal type_cast_2154_inst_req_1 : boolean;
  signal type_cast_2154_inst_ack_1 : boolean;
  signal SGT_f64_u1_2160_inst_req_0 : boolean;
  signal SGT_f64_u1_2160_inst_ack_0 : boolean;
  signal SGT_f64_u1_2160_inst_req_1 : boolean;
  signal SGT_f64_u1_2160_inst_ack_1 : boolean;
  signal if_stmt_2162_branch_req_0 : boolean;
  signal if_stmt_2162_branch_ack_1 : boolean;
  signal if_stmt_2162_branch_ack_0 : boolean;
  signal STORE_is_decoded_2169_store_0_req_0 : boolean;
  signal STORE_is_decoded_2169_store_0_ack_0 : boolean;
  signal STORE_is_decoded_2169_store_0_req_1 : boolean;
  signal STORE_is_decoded_2169_store_0_ack_1 : boolean;
  signal ptr_deref_2184_store_0_req_0 : boolean;
  signal ptr_deref_2184_store_0_ack_0 : boolean;
  signal ptr_deref_2184_store_0_req_1 : boolean;
  signal ptr_deref_2184_store_0_ack_1 : boolean;
  signal SLT_f64_u1_2194_inst_req_0 : boolean;
  signal SLT_f64_u1_2194_inst_ack_0 : boolean;
  signal SLT_f64_u1_2194_inst_req_1 : boolean;
  signal SLT_f64_u1_2194_inst_ack_1 : boolean;
  signal if_stmt_2196_branch_req_0 : boolean;
  signal if_stmt_2196_branch_ack_1 : boolean;
  signal if_stmt_2196_branch_ack_0 : boolean;
  signal ptr_deref_2205_load_0_req_0 : boolean;
  signal ptr_deref_2205_load_0_ack_0 : boolean;
  signal ptr_deref_2205_load_0_req_1 : boolean;
  signal ptr_deref_2205_load_0_ack_1 : boolean;
  signal ADD_u64_u64_2380_inst_req_1 : boolean;
  signal type_cast_2209_inst_req_0 : boolean;
  signal type_cast_2209_inst_ack_0 : boolean;
  signal type_cast_2209_inst_req_1 : boolean;
  signal type_cast_2209_inst_ack_1 : boolean;
  signal ADD_u64_u64_2394_inst_ack_0 : boolean;
  signal ADD_u64_u64_2394_inst_req_0 : boolean;
  signal addr_of_2385_final_reg_ack_1 : boolean;
  signal SLT_f64_u1_2215_inst_req_0 : boolean;
  signal SLT_f64_u1_2215_inst_ack_0 : boolean;
  signal addr_of_2385_final_reg_req_1 : boolean;
  signal SLT_f64_u1_2215_inst_req_1 : boolean;
  signal SLT_f64_u1_2215_inst_ack_1 : boolean;
  signal if_stmt_2217_branch_req_0 : boolean;
  signal addr_of_2385_final_reg_ack_0 : boolean;
  signal if_stmt_2217_branch_ack_1 : boolean;
  signal addr_of_2385_final_reg_req_0 : boolean;
  signal if_stmt_2217_branch_ack_0 : boolean;
  signal STORE_is_decoded_2224_store_0_req_0 : boolean;
  signal STORE_is_decoded_2224_store_0_ack_0 : boolean;
  signal STORE_is_decoded_2224_store_0_req_1 : boolean;
  signal STORE_is_decoded_2224_store_0_ack_1 : boolean;
  signal ADD_u64_u64_2365_inst_ack_1 : boolean;
  signal type_cast_2389_inst_ack_1 : boolean;
  signal type_cast_2389_inst_req_1 : boolean;
  signal type_cast_2250_inst_req_0 : boolean;
  signal ptr_deref_2239_store_0_req_0 : boolean;
  signal ptr_deref_2239_store_0_ack_0 : boolean;
  signal ptr_deref_2239_store_0_req_1 : boolean;
  signal ptr_deref_2239_store_0_ack_1 : boolean;
  signal type_cast_2252_inst_req_1 : boolean;
  signal ADD_u64_u64_2365_inst_req_1 : boolean;
  signal ADD_u64_u64_2258_inst_req_0 : boolean;
  signal ADD_u64_u64_2258_inst_ack_0 : boolean;
  signal ADD_u64_u64_2258_inst_req_1 : boolean;
  signal ADD_u64_u64_2258_inst_ack_1 : boolean;
  signal EQ_u64_u1_2263_inst_req_0 : boolean;
  signal EQ_u64_u1_2263_inst_ack_0 : boolean;
  signal EQ_u64_u1_2263_inst_req_1 : boolean;
  signal EQ_u64_u1_2263_inst_ack_1 : boolean;
  signal if_stmt_2265_branch_req_0 : boolean;
  signal if_stmt_2265_branch_ack_1 : boolean;
  signal if_stmt_2265_branch_ack_0 : boolean;
  signal if_stmt_2677_branch_ack_1 : boolean;
  signal EQ_u16_u1_2281_inst_req_0 : boolean;
  signal EQ_u16_u1_2281_inst_ack_0 : boolean;
  signal EQ_u16_u1_2281_inst_req_1 : boolean;
  signal EQ_u16_u1_2281_inst_ack_1 : boolean;
  signal if_stmt_2283_branch_req_0 : boolean;
  signal LOAD_Nitr_required_2685_load_0_req_0 : boolean;
  signal if_stmt_2283_branch_ack_1 : boolean;
  signal if_stmt_2283_branch_ack_0 : boolean;
  signal if_stmt_2677_branch_ack_0 : boolean;
  signal LOAD_Nitr_required_2685_load_0_ack_0 : boolean;
  signal LOAD_nrows_2291_load_0_req_0 : boolean;
  signal LOAD_nrows_2291_load_0_ack_0 : boolean;
  signal LOAD_nrows_2291_load_0_req_1 : boolean;
  signal LOAD_nrows_2291_load_0_ack_1 : boolean;
  signal EQ_u16_u1_2297_inst_req_0 : boolean;
  signal EQ_u16_u1_2297_inst_ack_0 : boolean;
  signal EQ_u16_u1_2297_inst_req_1 : boolean;
  signal EQ_u16_u1_2297_inst_ack_1 : boolean;
  signal LOAD_Nitr_required_2685_load_0_req_1 : boolean;
  signal LOAD_Nitr_required_2685_load_0_ack_1 : boolean;
  signal if_stmt_2299_branch_req_0 : boolean;
  signal if_stmt_2299_branch_ack_1 : boolean;
  signal if_stmt_2299_branch_ack_0 : boolean;
  signal type_cast_2308_inst_req_0 : boolean;
  signal type_cast_2308_inst_ack_0 : boolean;
  signal type_cast_2308_inst_req_1 : boolean;
  signal type_cast_2308_inst_ack_1 : boolean;
  signal ADD_u32_u32_2314_inst_req_0 : boolean;
  signal ADD_u32_u32_2314_inst_ack_0 : boolean;
  signal ADD_u32_u32_2314_inst_req_1 : boolean;
  signal ADD_u32_u32_2314_inst_ack_1 : boolean;
  signal UGT_u16_u1_2320_inst_req_0 : boolean;
  signal UGT_u16_u1_2320_inst_ack_0 : boolean;
  signal UGT_u16_u1_2320_inst_req_1 : boolean;
  signal UGT_u16_u1_2320_inst_ack_1 : boolean;
  signal ADD_u16_u16_2326_inst_req_0 : boolean;
  signal ADD_u16_u16_2326_inst_ack_0 : boolean;
  signal ADD_u16_u16_2326_inst_req_1 : boolean;
  signal ADD_u16_u16_2326_inst_ack_1 : boolean;
  signal type_cast_2330_inst_req_0 : boolean;
  signal type_cast_2330_inst_ack_0 : boolean;
  signal type_cast_2330_inst_req_1 : boolean;
  signal type_cast_2330_inst_ack_1 : boolean;
  signal ADD_u64_u64_2336_inst_req_0 : boolean;
  signal ADD_u64_u64_2336_inst_ack_0 : boolean;
  signal ADD_u64_u64_2336_inst_req_1 : boolean;
  signal ADD_u64_u64_2336_inst_ack_1 : boolean;
  signal MUX_2343_inst_req_0 : boolean;
  signal MUX_2343_inst_ack_0 : boolean;
  signal MUX_2343_inst_req_1 : boolean;
  signal MUX_2343_inst_ack_1 : boolean;
  signal ADD_u16_u16_2349_inst_req_0 : boolean;
  signal ADD_u16_u16_2349_inst_ack_0 : boolean;
  signal ADD_u16_u16_2349_inst_req_1 : boolean;
  signal ADD_u16_u16_2349_inst_ack_1 : boolean;
  signal type_cast_2353_inst_req_0 : boolean;
  signal type_cast_2353_inst_ack_0 : boolean;
  signal type_cast_2353_inst_req_1 : boolean;
  signal type_cast_2353_inst_ack_1 : boolean;
  signal ADD_u64_u64_2359_inst_req_0 : boolean;
  signal ADD_u64_u64_2359_inst_ack_0 : boolean;
  signal ADD_u64_u64_2359_inst_req_1 : boolean;
  signal ADD_u64_u64_2359_inst_ack_1 : boolean;
  signal ADD_u64_u64_2365_inst_req_0 : boolean;
  signal ADD_u64_u64_2365_inst_ack_0 : boolean;
  signal addr_of_2399_final_reg_req_0 : boolean;
  signal addr_of_2399_final_reg_ack_0 : boolean;
  signal addr_of_2399_final_reg_req_1 : boolean;
  signal addr_of_2399_final_reg_ack_1 : boolean;
  signal EQ_u32_u1_2404_inst_req_0 : boolean;
  signal EQ_u32_u1_2404_inst_ack_0 : boolean;
  signal EQ_u32_u1_2404_inst_req_1 : boolean;
  signal EQ_u32_u1_2404_inst_ack_1 : boolean;
  signal if_stmt_2406_branch_req_0 : boolean;
  signal if_stmt_2406_branch_ack_1 : boolean;
  signal if_stmt_2406_branch_ack_0 : boolean;
  signal ptr_deref_2415_load_0_req_0 : boolean;
  signal ptr_deref_2415_load_0_ack_0 : boolean;
  signal ptr_deref_2415_load_0_req_1 : boolean;
  signal ptr_deref_2415_load_0_ack_1 : boolean;
  signal SUB_u16_u16_2420_inst_req_0 : boolean;
  signal SUB_u16_u16_2420_inst_ack_0 : boolean;
  signal SUB_u16_u16_2420_inst_req_1 : boolean;
  signal SUB_u16_u16_2420_inst_ack_1 : boolean;
  signal ptr_deref_2426_load_0_req_0 : boolean;
  signal ptr_deref_2426_load_0_ack_0 : boolean;
  signal ptr_deref_2426_load_0_req_1 : boolean;
  signal ptr_deref_2426_load_0_ack_1 : boolean;
  signal ptr_deref_2430_load_0_req_0 : boolean;
  signal ptr_deref_2430_load_0_ack_0 : boolean;
  signal ptr_deref_2430_load_0_req_1 : boolean;
  signal ptr_deref_2430_load_0_ack_1 : boolean;
  signal SUB_u16_u16_2435_inst_req_0 : boolean;
  signal SUB_u16_u16_2435_inst_ack_0 : boolean;
  signal SUB_u16_u16_2435_inst_req_1 : boolean;
  signal SUB_u16_u16_2435_inst_ack_1 : boolean;
  signal EQ_u16_u1_2456_inst_req_0 : boolean;
  signal EQ_u16_u1_2456_inst_ack_0 : boolean;
  signal EQ_u16_u1_2456_inst_req_1 : boolean;
  signal EQ_u16_u1_2456_inst_ack_1 : boolean;
  signal if_stmt_2458_branch_req_0 : boolean;
  signal if_stmt_2458_branch_ack_1 : boolean;
  signal if_stmt_2458_branch_ack_0 : boolean;
  signal ADD_u16_u16_2469_inst_req_0 : boolean;
  signal ADD_u16_u16_2469_inst_ack_0 : boolean;
  signal ADD_u16_u16_2469_inst_req_1 : boolean;
  signal ADD_u16_u16_2469_inst_ack_1 : boolean;
  signal ADD_u16_u16_2484_inst_req_0 : boolean;
  signal ADD_u16_u16_2484_inst_ack_0 : boolean;
  signal ADD_u16_u16_2484_inst_req_1 : boolean;
  signal ADD_u16_u16_2484_inst_ack_1 : boolean;
  signal type_cast_2488_inst_req_0 : boolean;
  signal type_cast_2488_inst_ack_0 : boolean;
  signal type_cast_2488_inst_req_1 : boolean;
  signal type_cast_2488_inst_ack_1 : boolean;
  signal ADD_u64_u64_2494_inst_req_0 : boolean;
  signal ADD_u64_u64_2494_inst_ack_0 : boolean;
  signal ADD_u64_u64_2494_inst_req_1 : boolean;
  signal ADD_u64_u64_2494_inst_ack_1 : boolean;
  signal addr_of_2499_final_reg_req_0 : boolean;
  signal addr_of_2499_final_reg_ack_0 : boolean;
  signal addr_of_2499_final_reg_req_1 : boolean;
  signal addr_of_2499_final_reg_ack_1 : boolean;
  signal ptr_deref_2503_load_0_req_0 : boolean;
  signal ptr_deref_2503_load_0_ack_0 : boolean;
  signal ptr_deref_2503_load_0_req_1 : boolean;
  signal ptr_deref_2503_load_0_ack_1 : boolean;
  signal ADD_u16_u16_2509_inst_req_0 : boolean;
  signal ADD_u16_u16_2509_inst_ack_0 : boolean;
  signal ADD_u16_u16_2509_inst_req_1 : boolean;
  signal ADD_u16_u16_2509_inst_ack_1 : boolean;
  signal type_cast_2513_inst_req_0 : boolean;
  signal type_cast_2513_inst_ack_0 : boolean;
  signal type_cast_2513_inst_req_1 : boolean;
  signal type_cast_2513_inst_ack_1 : boolean;
  signal addr_of_2518_final_reg_req_0 : boolean;
  signal addr_of_2518_final_reg_ack_0 : boolean;
  signal addr_of_2518_final_reg_req_1 : boolean;
  signal addr_of_2518_final_reg_ack_1 : boolean;
  signal ptr_deref_2522_load_0_req_0 : boolean;
  signal ptr_deref_2522_load_0_ack_0 : boolean;
  signal ptr_deref_2522_load_0_req_1 : boolean;
  signal ptr_deref_2522_load_0_ack_1 : boolean;
  signal type_cast_2375_inst_req_0 : boolean;
  signal addr_of_2527_final_reg_req_0 : boolean;
  signal addr_of_2527_final_reg_ack_0 : boolean;
  signal addr_of_2527_final_reg_req_1 : boolean;
  signal addr_of_2527_final_reg_ack_1 : boolean;
  signal type_cast_2375_inst_ack_0 : boolean;
  signal type_cast_2250_inst_ack_1 : boolean;
  signal type_cast_2250_inst_req_1 : boolean;
  signal ptr_deref_2531_load_0_req_0 : boolean;
  signal ptr_deref_2531_load_0_ack_0 : boolean;
  signal phi_stmt_2369_req_0 : boolean;
  signal ptr_deref_2531_load_0_req_1 : boolean;
  signal ptr_deref_2531_load_0_ack_1 : boolean;
  signal type_cast_2375_inst_ack_1 : boolean;
  signal phi_stmt_2369_req_1 : boolean;
  signal SUB_f32_f32_2536_inst_req_0 : boolean;
  signal SUB_f32_f32_2536_inst_ack_0 : boolean;
  signal SUB_f32_f32_2536_inst_req_1 : boolean;
  signal SUB_f32_f32_2536_inst_ack_1 : boolean;
  signal phi_stmt_2245_req_1 : boolean;
  signal type_cast_2250_inst_ack_0 : boolean;
  signal type_cast_2252_inst_ack_1 : boolean;
  signal addr_of_2541_final_reg_req_0 : boolean;
  signal addr_of_2541_final_reg_ack_0 : boolean;
  signal addr_of_2541_final_reg_req_1 : boolean;
  signal addr_of_2541_final_reg_ack_1 : boolean;
  signal phi_stmt_2245_req_2 : boolean;
  signal ptr_deref_2544_store_0_req_0 : boolean;
  signal ptr_deref_2544_store_0_ack_0 : boolean;
  signal ptr_deref_2544_store_0_req_1 : boolean;
  signal ptr_deref_2544_store_0_ack_1 : boolean;
  signal ADD_u16_u16_2551_inst_req_0 : boolean;
  signal ADD_u16_u16_2551_inst_ack_0 : boolean;
  signal ADD_u16_u16_2551_inst_req_1 : boolean;
  signal ADD_u16_u16_2551_inst_ack_1 : boolean;
  signal EQ_u16_u1_2556_inst_req_0 : boolean;
  signal EQ_u16_u1_2556_inst_ack_0 : boolean;
  signal EQ_u16_u1_2556_inst_req_1 : boolean;
  signal EQ_u16_u1_2556_inst_ack_1 : boolean;
  signal if_stmt_2558_branch_req_0 : boolean;
  signal if_stmt_2558_branch_ack_1 : boolean;
  signal if_stmt_2558_branch_ack_0 : boolean;
  signal ADD_u64_u64_2571_inst_req_0 : boolean;
  signal ADD_u64_u64_2571_inst_ack_0 : boolean;
  signal ADD_u64_u64_2571_inst_req_1 : boolean;
  signal ADD_u64_u64_2571_inst_ack_1 : boolean;
  signal EQ_u64_u1_2576_inst_req_0 : boolean;
  signal EQ_u64_u1_2576_inst_ack_0 : boolean;
  signal EQ_u64_u1_2576_inst_req_1 : boolean;
  signal EQ_u64_u1_2576_inst_ack_1 : boolean;
  signal type_cast_2375_inst_req_1 : boolean;
  signal if_stmt_2578_branch_req_0 : boolean;
  signal if_stmt_2578_branch_ack_1 : boolean;
  signal if_stmt_2578_branch_ack_0 : boolean;
  signal ADD_u16_u16_2591_inst_req_0 : boolean;
  signal ADD_u16_u16_2591_inst_ack_0 : boolean;
  signal ADD_u16_u16_2591_inst_req_1 : boolean;
  signal ADD_u16_u16_2591_inst_ack_1 : boolean;
  signal STORE_Nitr_required_2608_store_0_req_0 : boolean;
  signal STORE_Nitr_required_2608_store_0_ack_0 : boolean;
  signal STORE_Nitr_required_2608_store_0_req_1 : boolean;
  signal STORE_Nitr_required_2608_store_0_ack_1 : boolean;
  signal EQ_u16_u1_2615_inst_req_0 : boolean;
  signal EQ_u16_u1_2615_inst_ack_0 : boolean;
  signal EQ_u16_u1_2615_inst_req_1 : boolean;
  signal EQ_u16_u1_2615_inst_ack_1 : boolean;
  signal if_stmt_2617_branch_req_0 : boolean;
  signal if_stmt_2617_branch_ack_1 : boolean;
  signal if_stmt_2617_branch_ack_0 : boolean;
  signal addr_of_2637_final_reg_req_0 : boolean;
  signal addr_of_2637_final_reg_ack_0 : boolean;
  signal addr_of_2637_final_reg_req_1 : boolean;
  signal addr_of_2637_final_reg_ack_1 : boolean;
  signal ADD_u64_u64_2643_inst_req_0 : boolean;
  signal ADD_u64_u64_2643_inst_ack_0 : boolean;
  signal ADD_u64_u64_2643_inst_req_1 : boolean;
  signal ADD_u64_u64_2643_inst_ack_1 : boolean;
  signal type_cast_2647_inst_req_0 : boolean;
  signal type_cast_2647_inst_ack_0 : boolean;
  signal type_cast_2647_inst_req_1 : boolean;
  signal type_cast_2647_inst_ack_1 : boolean;
  signal ADD_u64_u64_2653_inst_req_0 : boolean;
  signal ADD_u64_u64_2653_inst_ack_0 : boolean;
  signal ADD_u64_u64_2653_inst_req_1 : boolean;
  signal ADD_u64_u64_2653_inst_ack_1 : boolean;
  signal ptr_deref_2657_load_0_req_0 : boolean;
  signal ptr_deref_2657_load_0_ack_0 : boolean;
  signal ptr_deref_2657_load_0_req_1 : boolean;
  signal ptr_deref_2657_load_0_ack_1 : boolean;
  signal WPIPE_code_block_decoded_2659_inst_req_0 : boolean;
  signal WPIPE_code_block_decoded_2659_inst_ack_0 : boolean;
  signal WPIPE_code_block_decoded_2659_inst_req_1 : boolean;
  signal WPIPE_code_block_decoded_2659_inst_ack_1 : boolean;
  signal LOAD_ncols_2663_load_0_req_0 : boolean;
  signal LOAD_ncols_2663_load_0_ack_0 : boolean;
  signal LOAD_ncols_2663_load_0_req_1 : boolean;
  signal LOAD_ncols_2663_load_0_ack_1 : boolean;
  signal type_cast_2667_inst_req_0 : boolean;
  signal type_cast_2667_inst_ack_0 : boolean;
  signal type_cast_2667_inst_req_1 : boolean;
  signal type_cast_2667_inst_ack_1 : boolean;
  signal SLT_i32_u1_2675_inst_req_0 : boolean;
  signal SLT_i32_u1_2675_inst_ack_0 : boolean;
  signal SLT_i32_u1_2675_inst_req_1 : boolean;
  signal SLT_i32_u1_2675_inst_ack_1 : boolean;
  signal if_stmt_2677_branch_req_0 : boolean;
  signal WPIPE_nitr_required_2698_inst_req_0 : boolean;
  signal WPIPE_nitr_required_2698_inst_ack_0 : boolean;
  signal WPIPE_nitr_required_2698_inst_req_1 : boolean;
  signal WPIPE_nitr_required_2698_inst_ack_1 : boolean;
  signal phi_stmt_1375_req_0 : boolean;
  signal phi_stmt_1375_ack_0 : boolean;
  signal type_cast_1447_inst_req_0 : boolean;
  signal type_cast_1447_inst_ack_0 : boolean;
  signal type_cast_1447_inst_req_1 : boolean;
  signal type_cast_1447_inst_ack_1 : boolean;
  signal phi_stmt_1444_req_0 : boolean;
  signal phi_stmt_1444_ack_0 : boolean;
  signal type_cast_1510_inst_req_0 : boolean;
  signal type_cast_1510_inst_ack_0 : boolean;
  signal type_cast_1510_inst_req_1 : boolean;
  signal type_cast_1510_inst_ack_1 : boolean;
  signal phi_stmt_1504_req_1 : boolean;
  signal phi_stmt_1504_req_0 : boolean;
  signal phi_stmt_1504_ack_0 : boolean;
  signal phi_stmt_1561_req_0 : boolean;
  signal type_cast_1570_inst_req_0 : boolean;
  signal type_cast_1570_inst_ack_0 : boolean;
  signal type_cast_1570_inst_req_1 : boolean;
  signal type_cast_1570_inst_ack_1 : boolean;
  signal phi_stmt_1561_req_2 : boolean;
  signal phi_stmt_1561_req_1 : boolean;
  signal phi_stmt_1561_ack_0 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal phi_stmt_1619_req_1 : boolean;
  signal phi_stmt_1619_req_0 : boolean;
  signal phi_stmt_1619_ack_0 : boolean;
  signal type_cast_1693_inst_req_0 : boolean;
  signal type_cast_1693_inst_ack_0 : boolean;
  signal type_cast_1693_inst_req_1 : boolean;
  signal type_cast_1693_inst_ack_1 : boolean;
  signal phi_stmt_1690_req_0 : boolean;
  signal phi_stmt_1690_req_1 : boolean;
  signal phi_stmt_1690_ack_0 : boolean;
  signal phi_stmt_1700_req_0 : boolean;
  signal type_cast_1712_inst_req_0 : boolean;
  signal type_cast_1712_inst_ack_0 : boolean;
  signal type_cast_1712_inst_req_1 : boolean;
  signal type_cast_1712_inst_ack_1 : boolean;
  signal phi_stmt_1707_req_1 : boolean;
  signal type_cast_1718_inst_req_0 : boolean;
  signal type_cast_1718_inst_ack_0 : boolean;
  signal type_cast_1718_inst_req_1 : boolean;
  signal type_cast_1718_inst_ack_1 : boolean;
  signal phi_stmt_1713_req_1 : boolean;
  signal type_cast_1706_inst_req_0 : boolean;
  signal type_cast_1706_inst_ack_0 : boolean;
  signal type_cast_1706_inst_req_1 : boolean;
  signal type_cast_1706_inst_ack_1 : boolean;
  signal phi_stmt_1700_req_1 : boolean;
  signal type_cast_1710_inst_req_0 : boolean;
  signal type_cast_1710_inst_ack_0 : boolean;
  signal type_cast_1710_inst_req_1 : boolean;
  signal type_cast_1710_inst_ack_1 : boolean;
  signal phi_stmt_1707_req_0 : boolean;
  signal type_cast_1716_inst_req_0 : boolean;
  signal type_cast_1716_inst_ack_0 : boolean;
  signal type_cast_1716_inst_req_1 : boolean;
  signal type_cast_1716_inst_ack_1 : boolean;
  signal phi_stmt_1713_req_0 : boolean;
  signal phi_stmt_1700_ack_0 : boolean;
  signal phi_stmt_1707_ack_0 : boolean;
  signal phi_stmt_1713_ack_0 : boolean;
  signal type_cast_1791_inst_req_0 : boolean;
  signal type_cast_1791_inst_ack_0 : boolean;
  signal type_cast_1791_inst_req_1 : boolean;
  signal type_cast_1791_inst_ack_1 : boolean;
  signal phi_stmt_1785_req_1 : boolean;
  signal phi_stmt_1785_req_0 : boolean;
  signal phi_stmt_1785_ack_0 : boolean;
  signal type_cast_1881_inst_req_0 : boolean;
  signal type_cast_1881_inst_ack_0 : boolean;
  signal type_cast_1881_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_1 : boolean;
  signal phi_stmt_1875_req_1 : boolean;
  signal phi_stmt_1875_req_0 : boolean;
  signal phi_stmt_1875_ack_0 : boolean;
  signal type_cast_1967_inst_req_0 : boolean;
  signal type_cast_1967_inst_ack_0 : boolean;
  signal type_cast_1967_inst_req_1 : boolean;
  signal type_cast_1967_inst_ack_1 : boolean;
  signal phi_stmt_1961_req_1 : boolean;
  signal phi_stmt_1961_req_0 : boolean;
  signal phi_stmt_1961_ack_0 : boolean;
  signal type_cast_2252_inst_ack_0 : boolean;
  signal type_cast_2442_inst_req_0 : boolean;
  signal type_cast_2442_inst_ack_0 : boolean;
  signal type_cast_2252_inst_req_0 : boolean;
  signal type_cast_2064_inst_req_0 : boolean;
  signal type_cast_2064_inst_ack_0 : boolean;
  signal type_cast_2064_inst_req_1 : boolean;
  signal type_cast_2064_inst_ack_1 : boolean;
  signal phi_stmt_2061_req_0 : boolean;
  signal type_cast_2442_inst_req_1 : boolean;
  signal type_cast_2442_inst_ack_1 : boolean;
  signal phi_stmt_2061_ack_0 : boolean;
  signal phi_stmt_2272_ack_0 : boolean;
  signal type_cast_2115_inst_req_0 : boolean;
  signal type_cast_2115_inst_ack_0 : boolean;
  signal phi_stmt_2272_req_0 : boolean;
  signal type_cast_2115_inst_req_1 : boolean;
  signal type_cast_2115_inst_ack_1 : boolean;
  signal phi_stmt_2109_req_1 : boolean;
  signal type_cast_2275_inst_ack_1 : boolean;
  signal type_cast_2275_inst_req_1 : boolean;
  signal type_cast_2275_inst_ack_0 : boolean;
  signal type_cast_2108_inst_req_0 : boolean;
  signal type_cast_2108_inst_ack_0 : boolean;
  signal type_cast_2275_inst_req_0 : boolean;
  signal type_cast_2108_inst_req_1 : boolean;
  signal type_cast_2108_inst_ack_1 : boolean;
  signal phi_stmt_2102_req_1 : boolean;
  signal phi_stmt_2109_req_0 : boolean;
  signal phi_stmt_2102_req_0 : boolean;
  signal phi_stmt_2102_ack_0 : boolean;
  signal phi_stmt_2109_ack_0 : boolean;
  signal phi_stmt_2245_ack_0 : boolean;
  signal type_cast_2181_inst_req_0 : boolean;
  signal type_cast_2181_inst_ack_0 : boolean;
  signal type_cast_2181_inst_req_1 : boolean;
  signal type_cast_2181_inst_ack_1 : boolean;
  signal phi_stmt_2175_req_1 : boolean;
  signal phi_stmt_2245_req_0 : boolean;
  signal type_cast_2248_inst_ack_1 : boolean;
  signal phi_stmt_2175_req_0 : boolean;
  signal type_cast_2248_inst_req_1 : boolean;
  signal phi_stmt_2175_ack_0 : boolean;
  signal phi_stmt_2369_ack_0 : boolean;
  signal phi_stmt_2230_ack_0 : boolean;
  signal type_cast_2248_inst_ack_0 : boolean;
  signal type_cast_2248_inst_req_0 : boolean;
  signal type_cast_2236_inst_req_0 : boolean;
  signal type_cast_2236_inst_ack_0 : boolean;
  signal type_cast_2236_inst_req_1 : boolean;
  signal type_cast_2236_inst_ack_1 : boolean;
  signal phi_stmt_2230_req_1 : boolean;
  signal phi_stmt_2230_req_0 : boolean;
  signal phi_stmt_2439_req_0 : boolean;
  signal type_cast_2448_inst_req_0 : boolean;
  signal type_cast_2448_inst_ack_0 : boolean;
  signal type_cast_2448_inst_req_1 : boolean;
  signal type_cast_2448_inst_ack_1 : boolean;
  signal phi_stmt_2445_req_0 : boolean;
  signal type_cast_2444_inst_req_0 : boolean;
  signal type_cast_2444_inst_ack_0 : boolean;
  signal type_cast_2444_inst_req_1 : boolean;
  signal type_cast_2444_inst_ack_1 : boolean;
  signal phi_stmt_2439_req_1 : boolean;
  signal type_cast_2450_inst_req_0 : boolean;
  signal type_cast_2450_inst_ack_0 : boolean;
  signal type_cast_2450_inst_req_1 : boolean;
  signal type_cast_2450_inst_ack_1 : boolean;
  signal phi_stmt_2445_req_1 : boolean;
  signal phi_stmt_2439_ack_0 : boolean;
  signal phi_stmt_2445_ack_0 : boolean;
  signal type_cast_2479_inst_req_0 : boolean;
  signal type_cast_2479_inst_ack_0 : boolean;
  signal type_cast_2479_inst_req_1 : boolean;
  signal type_cast_2479_inst_ack_1 : boolean;
  signal phi_stmt_2473_req_1 : boolean;
  signal phi_stmt_2473_req_0 : boolean;
  signal phi_stmt_2473_ack_0 : boolean;
  signal type_cast_2598_inst_req_0 : boolean;
  signal type_cast_2598_inst_ack_0 : boolean;
  signal type_cast_2598_inst_req_1 : boolean;
  signal type_cast_2598_inst_ack_1 : boolean;
  signal phi_stmt_2595_req_0 : boolean;
  signal type_cast_2604_inst_req_0 : boolean;
  signal type_cast_2604_inst_ack_0 : boolean;
  signal type_cast_2604_inst_req_1 : boolean;
  signal type_cast_2604_inst_ack_1 : boolean;
  signal phi_stmt_2601_req_0 : boolean;
  signal type_cast_2600_inst_req_0 : boolean;
  signal type_cast_2600_inst_ack_0 : boolean;
  signal type_cast_2600_inst_req_1 : boolean;
  signal type_cast_2600_inst_ack_1 : boolean;
  signal phi_stmt_2595_req_1 : boolean;
  signal type_cast_2606_inst_req_0 : boolean;
  signal type_cast_2606_inst_ack_0 : boolean;
  signal type_cast_2606_inst_req_1 : boolean;
  signal type_cast_2606_inst_ack_1 : boolean;
  signal phi_stmt_2601_req_1 : boolean;
  signal phi_stmt_2595_ack_0 : boolean;
  signal phi_stmt_2601_ack_0 : boolean;
  signal type_cast_2629_inst_req_0 : boolean;
  signal type_cast_2629_inst_ack_0 : boolean;
  signal type_cast_2629_inst_req_1 : boolean;
  signal type_cast_2629_inst_ack_1 : boolean;
  signal phi_stmt_2626_req_0 : boolean;
  signal phi_stmt_2626_req_1 : boolean;
  signal phi_stmt_2626_ack_0 : boolean;
  signal type_cast_2696_inst_req_0 : boolean;
  signal type_cast_2696_inst_ack_0 : boolean;
  signal type_cast_2696_inst_req_1 : boolean;
  signal type_cast_2696_inst_ack_1 : boolean;
  signal phi_stmt_2689_req_2 : boolean;
  signal type_cast_2694_inst_req_0 : boolean;
  signal type_cast_2694_inst_ack_0 : boolean;
  signal type_cast_2694_inst_req_1 : boolean;
  signal type_cast_2694_inst_ack_1 : boolean;
  signal phi_stmt_2689_req_1 : boolean;
  signal type_cast_2692_inst_req_0 : boolean;
  signal type_cast_2692_inst_ack_0 : boolean;
  signal type_cast_2692_inst_req_1 : boolean;
  signal type_cast_2692_inst_ack_1 : boolean;
  signal phi_stmt_2689_req_0 : boolean;
  signal phi_stmt_2689_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "minSumDecode_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  minSumDecode_CP_6680_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "minSumDecode_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= minSumDecode_CP_6680_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= minSumDecode_CP_6680_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= minSumDecode_CP_6680_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  minSumDecode_CP_6680: Block -- control-path 
    signal minSumDecode_CP_6680_elements: BooleanArray(1231 downto 0);
    -- 
  begin -- 
    minSumDecode_CP_6680_elements(0) <= minSumDecode_CP_6680_start;
    minSumDecode_CP_6680_symbol <= minSumDecode_CP_6680_elements(1230);
    -- CP-element group 0:  transition  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (2) 
      -- CP-element group 0: 	 branch_block_stmt_1353/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	856 
    -- CP-element group 1:  members (2) 
      -- CP-element group 1: 	 branch_block_stmt_1353/bb_0_bb_1
      -- CP-element group 1: 	 branch_block_stmt_1353/branch_block_stmt_1353__entry__
      -- 
    minSumDecode_CP_6680_elements(1) <= minSumDecode_CP_6680_elements(0);
    -- CP-element group 2:  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	1230 
    -- CP-element group 2:  members (1) 
      -- CP-element group 2: 	 branch_block_stmt_1353/branch_block_stmt_1353__exit__
      -- 
    minSumDecode_CP_6680_elements(2) <= false; 
    -- CP-element group 3:  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	859 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	108 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_1353/call_stmt_1356__entry__
      -- CP-element group 3: 	 branch_block_stmt_1353/merge_stmt_1355__exit__
      -- 
    minSumDecode_CP_6680_elements(3) <= minSumDecode_CP_6680_elements(859);
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	110 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	111 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365__entry__
      -- CP-element group 4: 	 branch_block_stmt_1353/call_stmt_1356__exit__
      -- 
    minSumDecode_CP_6680_elements(4) <= minSumDecode_CP_6680_elements(110);
    -- CP-element group 5:  branch  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	115 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	116 
    -- CP-element group 5: 	117 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_1353/if_stmt_1366__entry__
      -- CP-element group 5: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365__exit__
      -- 
    minSumDecode_CP_6680_elements(5) <= minSumDecode_CP_6680_elements(115);
    -- CP-element group 6:  merge  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	862 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	863 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi
      -- CP-element group 6: 	 branch_block_stmt_1353/merge_stmt_1372__exit__
      -- 
    minSumDecode_CP_6680_elements(6) <= minSumDecode_CP_6680_elements(862);
    -- CP-element group 7:  place  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	868 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	125 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1353/do_while_stmt_1381__entry__
      -- CP-element group 7: 	 branch_block_stmt_1353/merge_stmt_1374__exit__
      -- 
    minSumDecode_CP_6680_elements(7) <= minSumDecode_CP_6680_elements(868);
    -- CP-element group 8:  branch  place  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	206 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	207 
    -- CP-element group 8: 	208 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_1353/if_stmt_1439__entry__
      -- CP-element group 8: 	 branch_block_stmt_1353/do_while_stmt_1381__exit__
      -- 
    minSumDecode_CP_6680_elements(8) <= minSumDecode_CP_6680_elements(206);
    -- CP-element group 9:  merge  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	213 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	869 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1353/merge_stmt_1443__entry__
      -- CP-element group 9: 	 branch_block_stmt_1353/if_stmt_1439__exit__
      -- 
    minSumDecode_CP_6680_elements(9) <= minSumDecode_CP_6680_elements(213);
    -- CP-element group 10:  merge  place  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	876 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	215 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_1353/assign_stmt_1454__entry__
      -- CP-element group 10: 	 branch_block_stmt_1353/merge_stmt_1443__exit__
      -- 
    minSumDecode_CP_6680_elements(10) <= minSumDecode_CP_6680_elements(876);
    -- CP-element group 11:  branch  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	217 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	218 
    -- CP-element group 11: 	219 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1353/if_stmt_1455__entry__
      -- CP-element group 11: 	 branch_block_stmt_1353/assign_stmt_1454__exit__
      -- 
    minSumDecode_CP_6680_elements(11) <= minSumDecode_CP_6680_elements(217);
    -- CP-element group 12:  merge  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	879 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	227 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501__entry__
      -- CP-element group 12: 	 branch_block_stmt_1353/merge_stmt_1461__exit__
      -- 
    minSumDecode_CP_6680_elements(12) <= minSumDecode_CP_6680_elements(879);
    -- CP-element group 13:  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	246 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	884 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501__exit__
      -- CP-element group 13: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6
      -- 
    minSumDecode_CP_6680_elements(13) <= minSumDecode_CP_6680_elements(246);
    -- CP-element group 14:  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	889 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	247 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551__entry__
      -- CP-element group 14: 	 branch_block_stmt_1353/merge_stmt_1503__exit__
      -- 
    minSumDecode_CP_6680_elements(14) <= minSumDecode_CP_6680_elements(889);
    -- CP-element group 15:  branch  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	265 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	266 
    -- CP-element group 15: 	267 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1353/if_stmt_1552__entry__
      -- CP-element group 15: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551__exit__
      -- 
    minSumDecode_CP_6680_elements(15) <= minSumDecode_CP_6680_elements(265);
    -- CP-element group 16:  merge  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	892 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	896 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit
      -- CP-element group 16: 	 branch_block_stmt_1353/merge_stmt_1558__exit__
      -- 
    minSumDecode_CP_6680_elements(16) <= minSumDecode_CP_6680_elements(892);
    -- CP-element group 17:  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	905 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	275 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580__entry__
      -- CP-element group 17: 	 branch_block_stmt_1353/merge_stmt_1560__exit__
      -- 
    minSumDecode_CP_6680_elements(17) <= minSumDecode_CP_6680_elements(905);
    -- CP-element group 18:  branch  place  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	279 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	280 
    -- CP-element group 18: 	281 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1353/if_stmt_1581__entry__
      -- CP-element group 18: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580__exit__
      -- 
    minSumDecode_CP_6680_elements(18) <= minSumDecode_CP_6680_elements(279);
    -- CP-element group 19:  merge  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	908 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	289 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1353/merge_stmt_1587__exit__
      -- CP-element group 19: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616__entry__
      -- 
    minSumDecode_CP_6680_elements(19) <= minSumDecode_CP_6680_elements(908);
    -- CP-element group 20:  place  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	301 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	913 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10
      -- CP-element group 20: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616__exit__
      -- 
    minSumDecode_CP_6680_elements(20) <= minSumDecode_CP_6680_elements(301);
    -- CP-element group 21:  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	918 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	302 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680__entry__
      -- CP-element group 21: 	 branch_block_stmt_1353/merge_stmt_1618__exit__
      -- 
    minSumDecode_CP_6680_elements(21) <= minSumDecode_CP_6680_elements(918);
    -- CP-element group 22:  branch  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	326 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	327 
    -- CP-element group 22: 	328 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680__exit__
      -- CP-element group 22: 	 branch_block_stmt_1353/if_stmt_1681__entry__
      -- 
    minSumDecode_CP_6680_elements(22) <= minSumDecode_CP_6680_elements(326);
    -- CP-element group 23:  merge  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	921 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	922 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader
      -- CP-element group 23: 	 branch_block_stmt_1353/merge_stmt_1687__exit__
      -- 
    minSumDecode_CP_6680_elements(23) <= minSumDecode_CP_6680_elements(921);
    -- CP-element group 24:  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	931 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	932 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit
      -- CP-element group 24: 	 branch_block_stmt_1353/merge_stmt_1689__exit__
      -- 
    minSumDecode_CP_6680_elements(24) <= minSumDecode_CP_6680_elements(931);
    -- CP-element group 25:  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	958 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	336 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733__entry__
      -- CP-element group 25: 	 branch_block_stmt_1353/merge_stmt_1699__exit__
      -- 
    minSumDecode_CP_6680_elements(25) <= minSumDecode_CP_6680_elements(958);
    -- CP-element group 26:  branch  place  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	343 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	344 
    -- CP-element group 26: 	345 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1353/if_stmt_1734__entry__
      -- CP-element group 26: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733__exit__
      -- 
    minSumDecode_CP_6680_elements(26) <= minSumDecode_CP_6680_elements(343);
    -- CP-element group 27:  merge  place  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	961 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	353 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1353/assign_stmt_1746__entry__
      -- CP-element group 27: 	 branch_block_stmt_1353/merge_stmt_1740__exit__
      -- 
    minSumDecode_CP_6680_elements(27) <= minSumDecode_CP_6680_elements(961);
    -- CP-element group 28:  branch  place  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	355 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	356 
    -- CP-element group 28: 	357 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1353/if_stmt_1747__entry__
      -- CP-element group 28: 	 branch_block_stmt_1353/assign_stmt_1746__exit__
      -- 
    minSumDecode_CP_6680_elements(28) <= minSumDecode_CP_6680_elements(355);
    -- CP-element group 29:  merge  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	964 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	365 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782__entry__
      -- CP-element group 29: 	 branch_block_stmt_1353/merge_stmt_1753__exit__
      -- 
    minSumDecode_CP_6680_elements(29) <= minSumDecode_CP_6680_elements(964);
    -- CP-element group 30:  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	377 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	969 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16
      -- CP-element group 30: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782__exit__
      -- 
    minSumDecode_CP_6680_elements(30) <= minSumDecode_CP_6680_elements(377);
    -- CP-element group 31:  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	974 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	378 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821__entry__
      -- CP-element group 31: 	 branch_block_stmt_1353/merge_stmt_1784__exit__
      -- 
    minSumDecode_CP_6680_elements(31) <= minSumDecode_CP_6680_elements(974);
    -- CP-element group 32:  branch  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	392 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	393 
    -- CP-element group 32: 	394 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1353/if_stmt_1822__entry__
      -- CP-element group 32: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821__exit__
      -- 
    minSumDecode_CP_6680_elements(32) <= minSumDecode_CP_6680_elements(392);
    -- CP-element group 33:  merge  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	977 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	979 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexitx_xloopexit_initialize_aPosteriorix_xexit
      -- CP-element group 33: 	 branch_block_stmt_1353/merge_stmt_1828__exit__
      -- 
    minSumDecode_CP_6680_elements(33) <= minSumDecode_CP_6680_elements(977);
    -- CP-element group 34:  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	981 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	402 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1353/assign_stmt_1836__entry__
      -- CP-element group 34: 	 branch_block_stmt_1353/merge_stmt_1830__exit__
      -- 
    minSumDecode_CP_6680_elements(34) <= minSumDecode_CP_6680_elements(981);
    -- CP-element group 35:  branch  place  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	404 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	405 
    -- CP-element group 35: 	406 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_1353/if_stmt_1837__entry__
      -- CP-element group 35: 	 branch_block_stmt_1353/assign_stmt_1836__exit__
      -- 
    minSumDecode_CP_6680_elements(35) <= minSumDecode_CP_6680_elements(404);
    -- CP-element group 36:  merge  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	984 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	414 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872__entry__
      -- CP-element group 36: 	 branch_block_stmt_1353/merge_stmt_1843__exit__
      -- 
    minSumDecode_CP_6680_elements(36) <= minSumDecode_CP_6680_elements(984);
    -- CP-element group 37:  place  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	426 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	989 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20
      -- CP-element group 37: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872__exit__
      -- 
    minSumDecode_CP_6680_elements(37) <= minSumDecode_CP_6680_elements(426);
    -- CP-element group 38:  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	994 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	427 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903__entry__
      -- CP-element group 38: 	 branch_block_stmt_1353/merge_stmt_1874__exit__
      -- 
    minSumDecode_CP_6680_elements(38) <= minSumDecode_CP_6680_elements(994);
    -- CP-element group 39:  branch  place  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	436 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	437 
    -- CP-element group 39: 	438 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903__exit__
      -- CP-element group 39: 	 branch_block_stmt_1353/if_stmt_1904__entry__
      -- 
    minSumDecode_CP_6680_elements(39) <= minSumDecode_CP_6680_elements(436);
    -- CP-element group 40:  merge  place  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	997 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	998 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexitx_xloopexit_initializeExtrinsicInfox_xexit
      -- CP-element group 40: 	 branch_block_stmt_1353/merge_stmt_1910__exit__
      -- 
    minSumDecode_CP_6680_elements(40) <= minSumDecode_CP_6680_elements(997);
    -- CP-element group 41:  place  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	1001 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	446 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1353/call_stmt_1913__entry__
      -- CP-element group 41: 	 branch_block_stmt_1353/merge_stmt_1912__exit__
      -- 
    minSumDecode_CP_6680_elements(41) <= minSumDecode_CP_6680_elements(1001);
    -- CP-element group 42:  place  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	448 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	449 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922__entry__
      -- CP-element group 42: 	 branch_block_stmt_1353/call_stmt_1913__exit__
      -- 
    minSumDecode_CP_6680_elements(42) <= minSumDecode_CP_6680_elements(448);
    -- CP-element group 43:  branch  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	453 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	454 
    -- CP-element group 43: 	455 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1353/if_stmt_1923__entry__
      -- CP-element group 43: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922__exit__
      -- 
    minSumDecode_CP_6680_elements(43) <= minSumDecode_CP_6680_elements(453);
    -- CP-element group 44:  merge  place  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	1004 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	463 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1353/merge_stmt_1929__exit__
      -- CP-element group 44: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958__entry__
      -- 
    minSumDecode_CP_6680_elements(44) <= minSumDecode_CP_6680_elements(1004);
    -- CP-element group 45:  place  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	475 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	1009 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24
      -- CP-element group 45: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958__exit__
      -- 
    minSumDecode_CP_6680_elements(45) <= minSumDecode_CP_6680_elements(475);
    -- CP-element group 46:  place  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	1014 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	476 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031__entry__
      -- CP-element group 46: 	 branch_block_stmt_1353/merge_stmt_1960__exit__
      -- 
    minSumDecode_CP_6680_elements(46) <= minSumDecode_CP_6680_elements(1014);
    -- CP-element group 47:  branch  place  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	506 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	507 
    -- CP-element group 47: 	508 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031__exit__
      -- CP-element group 47: 	 branch_block_stmt_1353/if_stmt_2032__entry__
      -- 
    minSumDecode_CP_6680_elements(47) <= minSumDecode_CP_6680_elements(506);
    -- CP-element group 48:  merge  place  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	1017 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	1019 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1353/merge_stmt_2038__exit__
      -- CP-element group 48: 	 branch_block_stmt_1353/update_aPosteriorix_xexitx_xloopexit_update_aPosteriorix_xexit
      -- 
    minSumDecode_CP_6680_elements(48) <= minSumDecode_CP_6680_elements(1017);
    -- CP-element group 49:  place  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	1021 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	516 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053__entry__
      -- CP-element group 49: 	 branch_block_stmt_1353/merge_stmt_2040__exit__
      -- 
    minSumDecode_CP_6680_elements(49) <= minSumDecode_CP_6680_elements(1021);
    -- CP-element group 50:  branch  place  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	523 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	524 
    -- CP-element group 50: 	525 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053__exit__
      -- CP-element group 50: 	 branch_block_stmt_1353/if_stmt_2054__entry__
      -- 
    minSumDecode_CP_6680_elements(50) <= minSumDecode_CP_6680_elements(523);
    -- CP-element group 51:  merge  place  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	1028 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	533 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1353/assign_stmt_2068__entry__
      -- CP-element group 51: 	 branch_block_stmt_1353/merge_stmt_2060__exit__
      -- 
    minSumDecode_CP_6680_elements(51) <= minSumDecode_CP_6680_elements(1028);
    -- CP-element group 52:  place  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	535 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	1219 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit
      -- CP-element group 52: 	 branch_block_stmt_1353/assign_stmt_2068__exit__
      -- 
    minSumDecode_CP_6680_elements(52) <= minSumDecode_CP_6680_elements(535);
    -- CP-element group 53:  place  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	1031 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	536 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099__entry__
      -- CP-element group 53: 	 branch_block_stmt_1353/merge_stmt_2070__exit__
      -- 
    minSumDecode_CP_6680_elements(53) <= minSumDecode_CP_6680_elements(1031);
    -- CP-element group 54:  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	548 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	1040 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29
      -- CP-element group 54: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099__exit__
      -- 
    minSumDecode_CP_6680_elements(54) <= minSumDecode_CP_6680_elements(548);
    -- CP-element group 55:  place  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	1050 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	549 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140__entry__
      -- CP-element group 55: 	 branch_block_stmt_1353/merge_stmt_2101__exit__
      -- 
    minSumDecode_CP_6680_elements(55) <= minSumDecode_CP_6680_elements(1050);
    -- CP-element group 56:  branch  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	560 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	561 
    -- CP-element group 56: 	562 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1353/if_stmt_2141__entry__
      -- CP-element group 56: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140__exit__
      -- 
    minSumDecode_CP_6680_elements(56) <= minSumDecode_CP_6680_elements(560);
    -- CP-element group 57:  merge  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	1053 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	570 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161__entry__
      -- CP-element group 57: 	 branch_block_stmt_1353/merge_stmt_2147__exit__
      -- 
    minSumDecode_CP_6680_elements(57) <= minSumDecode_CP_6680_elements(1053);
    -- CP-element group 58:  branch  place  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	576 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	577 
    -- CP-element group 58: 	578 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1353/if_stmt_2162__entry__
      -- CP-element group 58: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161__exit__
      -- 
    minSumDecode_CP_6680_elements(58) <= minSumDecode_CP_6680_elements(576);
    -- CP-element group 59:  merge  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	1056 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	586 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_1353/assign_stmt_2172__entry__
      -- CP-element group 59: 	 branch_block_stmt_1353/merge_stmt_2168__exit__
      -- 
    minSumDecode_CP_6680_elements(59) <= minSumDecode_CP_6680_elements(1056);
    -- CP-element group 60:  place  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	588 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	1061 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1353/assign_stmt_2172__exit__
      -- CP-element group 60: 	 branch_block_stmt_1353/bb_31_bb_32
      -- 
    minSumDecode_CP_6680_elements(60) <= minSumDecode_CP_6680_elements(588);
    -- CP-element group 61:  place  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	1066 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	589 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1353/assign_stmt_2187__entry__
      -- CP-element group 61: 	 branch_block_stmt_1353/merge_stmt_2174__exit__
      -- 
    minSumDecode_CP_6680_elements(61) <= minSumDecode_CP_6680_elements(1066);
    -- CP-element group 62:  place  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	591 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	1086 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1353/bb_32_bb_37
      -- CP-element group 62: 	 branch_block_stmt_1353/assign_stmt_2187__exit__
      -- 
    minSumDecode_CP_6680_elements(62) <= minSumDecode_CP_6680_elements(591);
    -- CP-element group 63:  place  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	1069 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	592 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1353/assign_stmt_2195__entry__
      -- CP-element group 63: 	 branch_block_stmt_1353/merge_stmt_2189__exit__
      -- 
    minSumDecode_CP_6680_elements(63) <= minSumDecode_CP_6680_elements(1069);
    -- CP-element group 64:  branch  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	594 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	595 
    -- CP-element group 64: 	596 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1353/if_stmt_2196__entry__
      -- CP-element group 64: 	 branch_block_stmt_1353/assign_stmt_2195__exit__
      -- 
    minSumDecode_CP_6680_elements(64) <= minSumDecode_CP_6680_elements(594);
    -- CP-element group 65:  merge  place  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	1072 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	604 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216__entry__
      -- CP-element group 65: 	 branch_block_stmt_1353/merge_stmt_2202__exit__
      -- 
    minSumDecode_CP_6680_elements(65) <= minSumDecode_CP_6680_elements(1072);
    -- CP-element group 66:  branch  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	610 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	611 
    -- CP-element group 66: 	612 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1353/if_stmt_2217__entry__
      -- CP-element group 66: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216__exit__
      -- 
    minSumDecode_CP_6680_elements(66) <= minSumDecode_CP_6680_elements(610);
    -- CP-element group 67:  merge  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	1075 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	620 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1353/assign_stmt_2227__entry__
      -- CP-element group 67: 	 branch_block_stmt_1353/merge_stmt_2223__exit__
      -- 
    minSumDecode_CP_6680_elements(67) <= minSumDecode_CP_6680_elements(1075);
    -- CP-element group 68:  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	622 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	1080 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1353/bb_35_bb_36
      -- CP-element group 68: 	 branch_block_stmt_1353/assign_stmt_2227__exit__
      -- 
    minSumDecode_CP_6680_elements(68) <= minSumDecode_CP_6680_elements(622);
    -- CP-element group 69:  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	1085 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	623 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1353/assign_stmt_2242__entry__
      -- CP-element group 69: 	 branch_block_stmt_1353/merge_stmt_2229__exit__
      -- 
    minSumDecode_CP_6680_elements(69) <= minSumDecode_CP_6680_elements(1085);
    -- CP-element group 70:  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	625 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	1094 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1353/bb_36_bb_37
      -- CP-element group 70: 	 branch_block_stmt_1353/assign_stmt_2242__exit__
      -- 
    minSumDecode_CP_6680_elements(70) <= minSumDecode_CP_6680_elements(625);
    -- CP-element group 71:  place  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	1100 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	626 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264__entry__
      -- CP-element group 71: 	 branch_block_stmt_1353/merge_stmt_2244__exit__
      -- 
    minSumDecode_CP_6680_elements(71) <= minSumDecode_CP_6680_elements(1100);
    -- CP-element group 72:  branch  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	630 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	631 
    -- CP-element group 72: 	632 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1353/if_stmt_2265__entry__
      -- CP-element group 72: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264__exit__
      -- 
    minSumDecode_CP_6680_elements(72) <= minSumDecode_CP_6680_elements(630);
    -- CP-element group 73:  merge  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	1107 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	640 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1353/assign_stmt_2282__entry__
      -- CP-element group 73: 	 branch_block_stmt_1353/merge_stmt_2271__exit__
      -- 
    minSumDecode_CP_6680_elements(73) <= minSumDecode_CP_6680_elements(1107);
    -- CP-element group 74:  branch  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	642 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	643 
    -- CP-element group 74: 	644 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1353/assign_stmt_2282__exit__
      -- CP-element group 74: 	 branch_block_stmt_1353/if_stmt_2283__entry__
      -- 
    minSumDecode_CP_6680_elements(74) <= minSumDecode_CP_6680_elements(642);
    -- CP-element group 75:  merge  place  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	1110 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	652 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298__entry__
      -- CP-element group 75: 	 branch_block_stmt_1353/merge_stmt_2289__exit__
      -- 
    minSumDecode_CP_6680_elements(75) <= minSumDecode_CP_6680_elements(1110);
    -- CP-element group 76:  branch  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	656 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	657 
    -- CP-element group 76: 	658 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1353/if_stmt_2299__entry__
      -- CP-element group 76: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298__exit__
      -- 
    minSumDecode_CP_6680_elements(76) <= minSumDecode_CP_6680_elements(656);
    -- CP-element group 77:  merge  place  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	1113 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	666 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366__entry__
      -- CP-element group 77: 	 branch_block_stmt_1353/merge_stmt_2305__exit__
      -- 
    minSumDecode_CP_6680_elements(77) <= minSumDecode_CP_6680_elements(1113);
    -- CP-element group 78:  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	690 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	1114 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366__exit__
      -- CP-element group 78: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41
      -- 
    minSumDecode_CP_6680_elements(78) <= minSumDecode_CP_6680_elements(690);
    -- CP-element group 79:  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	1123 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	691 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1353/merge_stmt_2368__exit__
      -- CP-element group 79: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405__entry__
      -- 
    minSumDecode_CP_6680_elements(79) <= minSumDecode_CP_6680_elements(1123);
    -- CP-element group 80:  branch  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	704 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	705 
    -- CP-element group 80: 	706 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405__exit__
      -- CP-element group 80: 	 branch_block_stmt_1353/if_stmt_2406__entry__
      -- 
    minSumDecode_CP_6680_elements(80) <= minSumDecode_CP_6680_elements(704);
    -- CP-element group 81:  merge  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	1126 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	714 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1353/merge_stmt_2412__exit__
      -- CP-element group 81: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421__entry__
      -- 
    minSumDecode_CP_6680_elements(81) <= minSumDecode_CP_6680_elements(1126);
    -- CP-element group 82:  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	718 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	1130 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421__exit__
      -- CP-element group 82: 	 branch_block_stmt_1353/bb_42_bb_44
      -- 
    minSumDecode_CP_6680_elements(82) <= minSumDecode_CP_6680_elements(718);
    -- CP-element group 83:  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1129 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	719 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1353/merge_stmt_2423__exit__
      -- CP-element group 83: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436__entry__
      -- 
    minSumDecode_CP_6680_elements(83) <= minSumDecode_CP_6680_elements(1129);
    -- CP-element group 84:  place  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	726 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	1138 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436__exit__
      -- CP-element group 84: 	 branch_block_stmt_1353/bb_43_bb_44
      -- 
    minSumDecode_CP_6680_elements(84) <= minSumDecode_CP_6680_elements(726);
    -- CP-element group 85:  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1150 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	727 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1353/merge_stmt_2438__exit__
      -- CP-element group 85: 	 branch_block_stmt_1353/assign_stmt_2457__entry__
      -- 
    minSumDecode_CP_6680_elements(85) <= minSumDecode_CP_6680_elements(1150);
    -- CP-element group 86:  branch  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	729 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	730 
    -- CP-element group 86: 	731 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1353/assign_stmt_2457__exit__
      -- CP-element group 86: 	 branch_block_stmt_1353/if_stmt_2458__entry__
      -- 
    minSumDecode_CP_6680_elements(86) <= minSumDecode_CP_6680_elements(729);
    -- CP-element group 87:  merge  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1153 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	739 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1353/merge_stmt_2464__exit__
      -- CP-element group 87: 	 branch_block_stmt_1353/assign_stmt_2470__entry__
      -- 
    minSumDecode_CP_6680_elements(87) <= minSumDecode_CP_6680_elements(1153);
    -- CP-element group 88:  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	741 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	1158 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1353/assign_stmt_2470__exit__
      -- CP-element group 88: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46
      -- 
    minSumDecode_CP_6680_elements(88) <= minSumDecode_CP_6680_elements(741);
    -- CP-element group 89:  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1163 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	742 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1353/merge_stmt_2472__exit__
      -- CP-element group 89: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557__entry__
      -- 
    minSumDecode_CP_6680_elements(89) <= minSumDecode_CP_6680_elements(1163);
    -- CP-element group 90:  branch  place  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	777 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	778 
    -- CP-element group 90: 	779 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557__exit__
      -- CP-element group 90: 	 branch_block_stmt_1353/if_stmt_2558__entry__
      -- 
    minSumDecode_CP_6680_elements(90) <= minSumDecode_CP_6680_elements(777);
    -- CP-element group 91:  merge  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1166 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	1168 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1353/merge_stmt_2564__exit__
      -- CP-element group 91: 	 branch_block_stmt_1353/xx_x_crit_edgex_xix_xloopexit_xx_x_crit_edgex_xi
      -- 
    minSumDecode_CP_6680_elements(91) <= minSumDecode_CP_6680_elements(1166);
    -- CP-element group 92:  place  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1170 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	787 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1353/merge_stmt_2566__exit__
      -- CP-element group 92: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577__entry__
      -- 
    minSumDecode_CP_6680_elements(92) <= minSumDecode_CP_6680_elements(1170);
    -- CP-element group 93:  branch  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	791 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	792 
    -- CP-element group 93: 	793 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577__exit__
      -- CP-element group 93: 	 branch_block_stmt_1353/if_stmt_2578__entry__
      -- 
    minSumDecode_CP_6680_elements(93) <= minSumDecode_CP_6680_elements(791);
    -- CP-element group 94:  merge  place  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1173 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	1175 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1353/merge_stmt_2584__exit__
      -- CP-element group 94: 	 branch_block_stmt_1353/updateMessagex_xexitx_xloopexit_updateMessagex_xexit
      -- 
    minSumDecode_CP_6680_elements(94) <= minSumDecode_CP_6680_elements(1173);
    -- CP-element group 95:  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1177 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	801 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1353/merge_stmt_2586__exit__
      -- CP-element group 95: 	 branch_block_stmt_1353/assign_stmt_2592__entry__
      -- 
    minSumDecode_CP_6680_elements(95) <= minSumDecode_CP_6680_elements(1177);
    -- CP-element group 96:  place  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	803 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	942 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1353/assign_stmt_2592__exit__
      -- CP-element group 96: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit
      -- 
    minSumDecode_CP_6680_elements(96) <= minSumDecode_CP_6680_elements(803);
    -- CP-element group 97:  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	1198 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	804 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1353/merge_stmt_2594__exit__
      -- CP-element group 97: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616__entry__
      -- 
    minSumDecode_CP_6680_elements(97) <= minSumDecode_CP_6680_elements(1198);
    -- CP-element group 98:  branch  place  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	809 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	810 
    -- CP-element group 98: 	811 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616__exit__
      -- CP-element group 98: 	 branch_block_stmt_1353/if_stmt_2617__entry__
      -- 
    minSumDecode_CP_6680_elements(98) <= minSumDecode_CP_6680_elements(809);
    -- CP-element group 99:  merge  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1201 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	1206 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1353/merge_stmt_2623__exit__
      -- CP-element group 99: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13
      -- 
    minSumDecode_CP_6680_elements(99) <= minSumDecode_CP_6680_elements(1201);
    -- CP-element group 100:  place  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1211 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	819 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_1353/merge_stmt_2625__exit__
      -- CP-element group 100: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658__entry__
      -- 
    minSumDecode_CP_6680_elements(100) <= minSumDecode_CP_6680_elements(1211);
    -- CP-element group 101:  place  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	830 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	831 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658__exit__
      -- CP-element group 101: 	 branch_block_stmt_1353/assign_stmt_2661__entry__
      -- 
    minSumDecode_CP_6680_elements(101) <= minSumDecode_CP_6680_elements(830);
    -- CP-element group 102:  place  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	833 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	834 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1353/assign_stmt_2661__exit__
      -- CP-element group 102: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676__entry__
      -- 
    minSumDecode_CP_6680_elements(102) <= minSumDecode_CP_6680_elements(833);
    -- CP-element group 103:  branch  place  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	840 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	841 
    -- CP-element group 103: 	842 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676__exit__
      -- CP-element group 103: 	 branch_block_stmt_1353/if_stmt_2677__entry__
      -- 
    minSumDecode_CP_6680_elements(103) <= minSumDecode_CP_6680_elements(840);
    -- CP-element group 104:  merge  place  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	1214 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	850 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1353/merge_stmt_2683__exit__
      -- CP-element group 104: 	 branch_block_stmt_1353/assign_stmt_2686__entry__
      -- 
    minSumDecode_CP_6680_elements(104) <= minSumDecode_CP_6680_elements(1214);
    -- CP-element group 105:  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	852 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	1223 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1353/assign_stmt_2686__exit__
      -- CP-element group 105: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit
      -- 
    minSumDecode_CP_6680_elements(105) <= minSumDecode_CP_6680_elements(852);
    -- CP-element group 106:  place  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1229 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	853 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1353/merge_stmt_2688__exit__
      -- CP-element group 106: 	 branch_block_stmt_1353/assign_stmt_2700__entry__
      -- 
    minSumDecode_CP_6680_elements(106) <= minSumDecode_CP_6680_elements(1229);
    -- CP-element group 107:  place  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	855 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	857 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1353/assign_stmt_2700__exit__
      -- CP-element group 107: 	 branch_block_stmt_1353/send_outputx_xexit_bb_1
      -- 
    minSumDecode_CP_6680_elements(107) <= minSumDecode_CP_6680_elements(855);
    -- CP-element group 108:  fork  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	3 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (7) 
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/$entry
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_update_start_
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Sample/crr
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Update/ccr
      -- 
    crr_6961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(108), ack => call_stmt_1356_call_req_0); -- 
    ccr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(108), ack => call_stmt_1356_call_req_1); -- 
    minSumDecode_CP_6680_elements(108) <= minSumDecode_CP_6680_elements(3);
    -- CP-element group 109:  transition  input  no-bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Sample/cra
      -- 
    cra_6962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1356_call_ack_0, ack => minSumDecode_CP_6680_elements(109)); -- 
    -- CP-element group 110:  transition  input  no-bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	4 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_1353/call_stmt_1356/$exit
      -- CP-element group 110: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1353/call_stmt_1356/call_stmt_1356_Update/cca
      -- 
    cca_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1356_call_ack_1, ack => minSumDecode_CP_6680_elements(110)); -- 
    -- CP-element group 111:  fork  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	4 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	115 
    -- CP-element group 111:  members (16) 
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_word_address_calculated
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_root_address_calculated
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/word_0/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/word_0/rr
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/word_0/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/word_0/cr
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Update/cr
      -- 
    cr_6997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(111), ack => LOAD_ncols_1358_load_0_req_1); -- 
    rr_6986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(111), ack => LOAD_ncols_1358_load_0_req_0); -- 
    cr_7016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(111), ack => EQ_u16_u1_1364_inst_req_1); -- 
    minSumDecode_CP_6680_elements(111) <= minSumDecode_CP_6680_elements(4);
    -- CP-element group 112:  transition  input  no-bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Sample/word_access_start/word_0/ra
      -- 
    ra_6987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_1358_load_0_ack_0, ack => minSumDecode_CP_6680_elements(112)); -- 
    -- CP-element group 113:  transition  input  output  no-bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (12) 
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/$exit
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/LOAD_ncols_1358_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/LOAD_ncols_1358_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/LOAD_ncols_1358_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/LOAD_ncols_1358_Update/LOAD_ncols_1358_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Sample/rr
      -- 
    ca_6998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_1358_load_0_ack_1, ack => minSumDecode_CP_6680_elements(113)); -- 
    rr_7011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(113), ack => EQ_u16_u1_1364_inst_req_0); -- 
    -- CP-element group 114:  transition  input  no-bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Sample/ra
      -- 
    ra_7012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1364_inst_ack_0, ack => minSumDecode_CP_6680_elements(114)); -- 
    -- CP-element group 115:  transition  input  no-bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	111 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	5 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/$exit
      -- CP-element group 115: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1353/assign_stmt_1359_to_assign_stmt_1365/EQ_u16_u1_1364_Update/ca
      -- 
    ca_7017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1364_inst_ack_1, ack => minSumDecode_CP_6680_elements(115)); -- 
    -- CP-element group 116:  transition  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	5 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1353/if_stmt_1366_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(116) <= minSumDecode_CP_6680_elements(5);
    -- CP-element group 117:  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	5 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1353/if_stmt_1366_eval_test/$entry
      -- CP-element group 117: 	 branch_block_stmt_1353/if_stmt_1366_eval_test/$exit
      -- CP-element group 117: 	 branch_block_stmt_1353/if_stmt_1366_eval_test/branch_req
      -- 
    branch_req_7025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(117), ack => if_stmt_1366_branch_req_0); -- 
    minSumDecode_CP_6680_elements(117) <= minSumDecode_CP_6680_elements(5);
    -- CP-element group 118:  branch  place  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	121 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1353/R_iNsTr_3_1367_place
      -- 
    minSumDecode_CP_6680_elements(118) <= minSumDecode_CP_6680_elements(117);
    -- CP-element group 119:  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1353/if_stmt_1366_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(119) <= minSumDecode_CP_6680_elements(118);
    -- CP-element group 120:  transition  input  no-bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1353/if_stmt_1366_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_1353/if_stmt_1366_if_link/if_choice_transition
      -- 
    if_choice_transition_7030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1366_branch_ack_1, ack => minSumDecode_CP_6680_elements(120)); -- 
    -- CP-element group 121:  transition  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	118 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1353/if_stmt_1366_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(121) <= minSumDecode_CP_6680_elements(118);
    -- CP-element group 122:  transition  input  no-bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1353/if_stmt_1366_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_1353/if_stmt_1366_else_link/else_choice_transition
      -- 
    else_choice_transition_7034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1366_branch_ack_0, ack => minSumDecode_CP_6680_elements(122)); -- 
    -- CP-element group 123:  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	893 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit
      -- 
    minSumDecode_CP_6680_elements(123) <= minSumDecode_CP_6680_elements(120);
    -- CP-element group 124:  place  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	860 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1353/bb_1_bbx_xnphx_xix_xpreheader
      -- 
    minSumDecode_CP_6680_elements(124) <= minSumDecode_CP_6680_elements(122);
    -- CP-element group 125:  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	7 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1353/do_while_stmt_1381/$entry
      -- 
    minSumDecode_CP_6680_elements(125) <= minSumDecode_CP_6680_elements(7);
    -- CP-element group 126:  place  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	132 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381__entry__
      -- 
    minSumDecode_CP_6680_elements(126) <= minSumDecode_CP_6680_elements(125);
    -- CP-element group 127:  merge  place  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	206 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381__exit__
      -- 
    -- Element group minSumDecode_CP_6680_elements(127) is bound as output of CP function.
    -- CP-element group 128:  merge  place  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_back
      -- 
    -- Element group minSumDecode_CP_6680_elements(128) is bound as output of CP function.
    -- CP-element group 129:  branch  place  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	134 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	202 
    -- CP-element group 129: 	204 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1353/do_while_stmt_1381/condition_done
      -- 
    minSumDecode_CP_6680_elements(129) <= minSumDecode_CP_6680_elements(134);
    -- CP-element group 130:  branch  place  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	1231 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_body_done
      -- 
    minSumDecode_CP_6680_elements(130) <= minSumDecode_CP_6680_elements(1231);
    -- CP-element group 131:  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	140 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/back_edge_to_loop_body
      -- 
    minSumDecode_CP_6680_elements(131) <= minSumDecode_CP_6680_elements(128);
    -- CP-element group 132:  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	126 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	142 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/first_time_through_loop_body
      -- 
    minSumDecode_CP_6680_elements(132) <= minSumDecode_CP_6680_elements(126);
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	136 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	159 
    -- CP-element group 133: 	166 
    -- CP-element group 133: 	171 
    -- CP-element group 133: 	175 
    -- CP-element group 133: 	179 
    -- CP-element group 133: 	183 
    -- CP-element group 133: 	186 
    -- CP-element group 133: 	187 
    -- CP-element group 133: 	191 
    -- CP-element group 133: 	195 
    -- CP-element group 133: 	199 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/$entry
      -- CP-element group 133: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/loop_body_start
      -- CP-element group 133: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_root_address_calculated
      -- 
    -- Element group minSumDecode_CP_6680_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	137 
    -- CP-element group 134: 	197 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	129 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/condition_evaluated
      -- 
    condition_evaluated_7051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(134), ack => do_while_stmt_1381_branch_req_0); -- 
    minSumDecode_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 16);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(137) & minSumDecode_CP_6680_elements(197);
      gj_minSumDecode_cp_element_group_134 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/aggregated_phi_sample_req
      -- CP-element group 135: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_sample_start__ps
      -- 
    minSumDecode_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(136) & minSumDecode_CP_6680_elements(139);
      gj_minSumDecode_cp_element_group_135 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  no-bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	133 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: 	165 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_sample_start_
      -- 
    minSumDecode_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(138) & minSumDecode_CP_6680_elements(165);
      gj_minSumDecode_cp_element_group_136 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  fork  transition  no-bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	133 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	160 
    -- CP-element group 137: 	164 
    -- CP-element group 137: 	172 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	134 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/aggregated_phi_update_req
      -- CP-element group 137: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_update_start__ps
      -- 
    minSumDecode_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 16,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 1,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(139) & minSumDecode_CP_6680_elements(160) & minSumDecode_CP_6680_elements(164) & minSumDecode_CP_6680_elements(172);
      gj_minSumDecode_cp_element_group_137 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	163 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/aggregated_phi_sample_ack
      -- CP-element group 138: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_sample_completed__ps
      -- 
    -- Element group minSumDecode_CP_6680_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	158 
    -- CP-element group 139: 	162 
    -- CP-element group 139: 	170 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/aggregated_phi_update_ack
      -- CP-element group 139: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_update_completed__ps
      -- 
    -- Element group minSumDecode_CP_6680_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	131 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_loopback_trigger
      -- 
    minSumDecode_CP_6680_elements(140) <= minSumDecode_CP_6680_elements(131);
    -- CP-element group 141:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_loopback_sample_req
      -- 
    phi_stmt_1383_loopback_sample_req_7066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1383_loopback_sample_req_7066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(141), ack => phi_stmt_1383_req_0); -- 
    -- Element group minSumDecode_CP_6680_elements(141) is bound as output of CP function.
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	132 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_entry_trigger
      -- 
    minSumDecode_CP_6680_elements(142) <= minSumDecode_CP_6680_elements(132);
    -- CP-element group 143:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_entry_sample_req
      -- 
    phi_stmt_1383_entry_sample_req_7068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1383_entry_sample_req_7068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(143), ack => phi_stmt_1383_req_1); -- 
    -- Element group minSumDecode_CP_6680_elements(143) is bound as output of CP function.
    -- CP-element group 144:  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_merged_reqs
      -- 
    -- Element group minSumDecode_CP_6680_elements(144) is bound as output of CP function.
    -- CP-element group 145:  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_entry_sample_req__merge_in
      -- 
    minSumDecode_CP_6680_elements(145) <= minSumDecode_CP_6680_elements(143);
    -- CP-element group 146:  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_loopback_sample_req__merge_in
      -- 
    minSumDecode_CP_6680_elements(146) <= minSumDecode_CP_6680_elements(141);
    -- CP-element group 147:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	1231 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_phi_mux_ack
      -- 
    phi_stmt_1383_phi_mux_ack_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1383_ack_0, ack => minSumDecode_CP_6680_elements(147)); -- 
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_sample_start__ps
      -- 
    -- Element group minSumDecode_CP_6680_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_update_start__ps
      -- 
    -- Element group minSumDecode_CP_6680_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Sample/rr
      -- 
    rr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(150), ack => type_cast_1386_inst_req_0); -- 
    minSumDecode_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(148) & minSumDecode_CP_6680_elements(152);
      gj_minSumDecode_cp_element_group_150 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Update/cr
      -- 
    cr_7091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(151), ack => type_cast_1386_inst_req_1); -- 
    minSumDecode_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(149) & minSumDecode_CP_6680_elements(153);
      gj_minSumDecode_cp_element_group_151 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Sample/ra
      -- 
    ra_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => minSumDecode_CP_6680_elements(152)); -- 
    -- CP-element group 153:  join  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1386_Update/ca
      -- 
    ca_7092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => minSumDecode_CP_6680_elements(153)); -- 
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_sample_start__ps
      -- CP-element group 154: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Sample/req
      -- 
    req_7104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(154), ack => iNsTr_13_at_entry_1375_1387_buf_req_0); -- 
    -- Element group minSumDecode_CP_6680_elements(154) is bound as output of CP function.
    -- CP-element group 155:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_update_start__ps
      -- CP-element group 155: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Update/req
      -- 
    req_7109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(155), ack => iNsTr_13_at_entry_1375_1387_buf_req_1); -- 
    -- Element group minSumDecode_CP_6680_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (4) 
      -- CP-element group 156: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_sample_completed__ps
      -- CP-element group 156: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Sample/ack
      -- 
    ack_7105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iNsTr_13_at_entry_1375_1387_buf_ack_0, ack => minSumDecode_CP_6680_elements(156)); -- 
    -- CP-element group 157:  join  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_update_completed__ps
      -- CP-element group 157: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/R_iNsTr_13_at_entry_1387_Update/ack
      -- 
    ack_7110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iNsTr_13_at_entry_1375_1387_buf_ack_1, ack => minSumDecode_CP_6680_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	139 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Sample/rr
      -- 
    rr_7119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(158), ack => ADD_u8_u8_1393_inst_req_0); -- 
    minSumDecode_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(139) & minSumDecode_CP_6680_elements(160);
      gj_minSumDecode_cp_element_group_158 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	133 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	184 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Update/cr
      -- 
    cr_7124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(159), ack => ADD_u8_u8_1393_inst_req_1); -- 
    minSumDecode_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(161) & minSumDecode_CP_6680_elements(184);
      gj_minSumDecode_cp_element_group_159 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	137 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Sample/ra
      -- 
    ra_7120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_1393_inst_ack_0, ack => minSumDecode_CP_6680_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	182 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1393_Update/ca
      -- 
    ca_7125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_1393_inst_ack_1, ack => minSumDecode_CP_6680_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	139 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Sample/rr
      -- 
    rr_7133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(162), ack => ADD_u8_u8_1399_inst_req_0); -- 
    minSumDecode_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(139) & minSumDecode_CP_6680_elements(164);
      gj_minSumDecode_cp_element_group_162 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	138 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Update/cr
      -- 
    cr_7138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(163), ack => ADD_u8_u8_1399_inst_req_1); -- 
    minSumDecode_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(138) & minSumDecode_CP_6680_elements(165);
      gj_minSumDecode_cp_element_group_163 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	137 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Sample/ra
      -- 
    ra_7134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_1399_inst_ack_0, ack => minSumDecode_CP_6680_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	1231 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	136 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ADD_u8_u8_1399_Update/ca
      -- 
    ca_7139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_1399_inst_ack_1, ack => minSumDecode_CP_6680_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	133 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Sample/rr
      -- 
    rr_7147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(166), ack => RPIPE_code_block_in_1402_inst_req_0); -- 
    minSumDecode_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(168);
      gj_minSumDecode_cp_element_group_166 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: 	180 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_update_start_
      -- CP-element group 167: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Update/cr
      -- 
    cr_7152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(167), ack => RPIPE_code_block_in_1402_inst_req_1); -- 
    minSumDecode_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(168) & minSumDecode_CP_6680_elements(169) & minSumDecode_CP_6680_elements(180);
      gj_minSumDecode_cp_element_group_167 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Sample/ra
      -- 
    ra_7148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_code_block_in_1402_inst_ack_0, ack => minSumDecode_CP_6680_elements(168)); -- 
    -- CP-element group 169:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	178 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/RPIPE_code_block_in_1402_Update/ca
      -- 
    ca_7153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_code_block_in_1402_inst_ack_1, ack => minSumDecode_CP_6680_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	139 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Sample/rr
      -- 
    rr_7161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(170), ack => type_cast_1406_inst_req_0); -- 
    minSumDecode_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(139) & minSumDecode_CP_6680_elements(172);
      gj_minSumDecode_cp_element_group_170 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	133 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Update/cr
      -- 
    cr_7166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(171), ack => type_cast_1406_inst_req_1); -- 
    minSumDecode_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(173);
      gj_minSumDecode_cp_element_group_171 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	137 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Sample/ra
      -- 
    ra_7162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => minSumDecode_CP_6680_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (24) 
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1406_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_offset_calculated
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_resized_0
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_scaled_0
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_computed_0
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_resize_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_resize_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_resize_0/index_resize_req
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_resize_0/index_resize_ack
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_scale_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_scale_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_scale_0/scale_rename_req
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_index_scale_0/scale_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_final_index_sum_regn/$entry
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_final_index_sum_regn/$exit
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_final_index_sum_regn/req
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_final_index_sum_regn/ack
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/array_obj_ref_1410_base_plus_offset/sum_rename_ack
      -- 
    ca_7167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => minSumDecode_CP_6680_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_request/$entry
      -- CP-element group 174: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_request/req
      -- 
    req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(174), ack => addr_of_1411_final_reg_req_0); -- 
    minSumDecode_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(173) & minSumDecode_CP_6680_elements(176);
      gj_minSumDecode_cp_element_group_174 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	133 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	180 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_complete/$entry
      -- CP-element group 175: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_complete/req
      -- 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(175), ack => addr_of_1411_final_reg_req_1); -- 
    minSumDecode_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(177) & minSumDecode_CP_6680_elements(180);
      gj_minSumDecode_cp_element_group_175 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	1231 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_request/$exit
      -- CP-element group 176: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_request/ack
      -- 
    ack_7201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1411_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (19) 
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_complete/$exit
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/addr_of_1411_complete/ack
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_word_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_root_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_address_resized
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_addr_resize/$entry
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_addr_resize/$exit
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_addr_resize/base_resize_req
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_addr_resize/base_resize_ack
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_plus_offset/$entry
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_plus_offset/$exit
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_plus_offset/sum_rename_req
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_base_plus_offset/sum_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_word_addrgen/$entry
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_word_addrgen/$exit
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_word_addrgen/root_register_req
      -- CP-element group 177: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_word_addrgen/root_register_ack
      -- 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1411_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	169 
    -- CP-element group 178: 	177 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/ptr_deref_1414_Split/$entry
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/ptr_deref_1414_Split/$exit
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/ptr_deref_1414_Split/split_req
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/ptr_deref_1414_Split/split_ack
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/$entry
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/word_0/$entry
      -- CP-element group 178: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/word_0/rr
      -- 
    rr_7244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(178), ack => ptr_deref_1414_store_0_req_0); -- 
    minSumDecode_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 16,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(169) & minSumDecode_CP_6680_elements(177) & minSumDecode_CP_6680_elements(180);
      gj_minSumDecode_cp_element_group_178 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	133 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (5) 
      -- CP-element group 179: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/$entry
      -- CP-element group 179: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/word_0/$entry
      -- CP-element group 179: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/word_0/cr
      -- 
    cr_7255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(179), ack => ptr_deref_1414_store_0_req_1); -- 
    minSumDecode_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(181);
      gj_minSumDecode_cp_element_group_179 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	167 
    -- CP-element group 180: 	175 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/$exit
      -- CP-element group 180: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/word_0/$exit
      -- CP-element group 180: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Sample/word_access_start/word_0/ra
      -- 
    ra_7245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_store_0_ack_0, ack => minSumDecode_CP_6680_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	1231 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ptr_deref_1414_Update/word_access_complete/word_0/ca
      -- 
    ca_7256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_store_0_ack_1, ack => minSumDecode_CP_6680_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	161 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Sample/rr
      -- 
    rr_7264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(182), ack => type_cast_1419_inst_req_0); -- 
    minSumDecode_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(161) & minSumDecode_CP_6680_elements(184);
      gj_minSumDecode_cp_element_group_182 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	133 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	196 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Update/cr
      -- 
    cr_7269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(183), ack => type_cast_1419_inst_req_1); -- 
    minSumDecode_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(185) & minSumDecode_CP_6680_elements(196);
      gj_minSumDecode_cp_element_group_183 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	159 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Sample/ra
      -- 
    ra_7265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_0, ack => minSumDecode_CP_6680_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	194 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1419_Update/ca
      -- 
    ca_7270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_1, ack => minSumDecode_CP_6680_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	133 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/$entry
      -- CP-element group 186: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/word_0/$entry
      -- CP-element group 186: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/word_0/rr
      -- 
    rr_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(186), ack => LOAD_ncols_1422_load_0_req_0); -- 
    minSumDecode_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(188);
      gj_minSumDecode_cp_element_group_186 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	133 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: 	192 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (5) 
      -- CP-element group 187: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/$entry
      -- CP-element group 187: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/word_0/$entry
      -- CP-element group 187: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/word_0/cr
      -- 
    cr_7297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(187), ack => LOAD_ncols_1422_load_0_req_1); -- 
    minSumDecode_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(189) & minSumDecode_CP_6680_elements(192);
      gj_minSumDecode_cp_element_group_187 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (5) 
      -- CP-element group 188: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/$exit
      -- CP-element group 188: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/word_0/$exit
      -- CP-element group 188: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Sample/word_access_start/word_0/ra
      -- 
    ra_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_1422_load_0_ack_0, ack => minSumDecode_CP_6680_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (9) 
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/$exit
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/word_0/$exit
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/word_access_complete/word_0/ca
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/LOAD_ncols_1422_Merge/$entry
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/LOAD_ncols_1422_Merge/$exit
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/LOAD_ncols_1422_Merge/merge_req
      -- CP-element group 189: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/LOAD_ncols_1422_Update/LOAD_ncols_1422_Merge/merge_ack
      -- 
    ca_7298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_1422_load_0_ack_1, ack => minSumDecode_CP_6680_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Sample/rr
      -- 
    rr_7311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(190), ack => type_cast_1426_inst_req_0); -- 
    minSumDecode_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(189) & minSumDecode_CP_6680_elements(192);
      gj_minSumDecode_cp_element_group_190 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	133 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: 	196 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_update_start_
      -- CP-element group 191: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Update/cr
      -- 
    cr_7316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(191), ack => type_cast_1426_inst_req_1); -- 
    minSumDecode_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(193) & minSumDecode_CP_6680_elements(196);
      gj_minSumDecode_cp_element_group_191 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	187 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Sample/ra
      -- 
    ra_7312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_0, ack => minSumDecode_CP_6680_elements(192)); -- 
    -- CP-element group 193:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/type_cast_1426_Update/ca
      -- 
    ca_7317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_1, ack => minSumDecode_CP_6680_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	185 
    -- CP-element group 194: 	193 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Sample/rr
      -- 
    rr_7325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(194), ack => ULT_u32_u1_1431_inst_req_0); -- 
    minSumDecode_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 16,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(185) & minSumDecode_CP_6680_elements(193) & minSumDecode_CP_6680_elements(196);
      gj_minSumDecode_cp_element_group_194 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	133 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: 	200 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Update/cr
      -- 
    cr_7330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(195), ack => ULT_u32_u1_1431_inst_req_1); -- 
    minSumDecode_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 16,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(197) & minSumDecode_CP_6680_elements(200);
      gj_minSumDecode_cp_element_group_195 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	183 
    -- CP-element group 196: 	191 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Sample/ra
      -- 
    ra_7326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_1431_inst_ack_0, ack => minSumDecode_CP_6680_elements(196)); -- 
    -- CP-element group 197:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	134 
    -- CP-element group 197: 	198 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/ULT_u32_u1_1431_Update/ca
      -- 
    ca_7331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u32_u1_1431_inst_ack_1, ack => minSumDecode_CP_6680_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Sample/rr
      -- 
    rr_7339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(198), ack => NOT_u1_u1_1435_inst_req_0); -- 
    minSumDecode_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(197) & minSumDecode_CP_6680_elements(200);
      gj_minSumDecode_cp_element_group_198 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  no-bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	133 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	201 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_update_start_
      -- CP-element group 199: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Update/cr
      -- 
    cr_7344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(199), ack => NOT_u1_u1_1435_inst_req_1); -- 
    minSumDecode_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 16,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(133) & minSumDecode_CP_6680_elements(201);
      gj_minSumDecode_cp_element_group_199 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Sample/ra
      -- 
    ra_7340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1435_inst_ack_0, ack => minSumDecode_CP_6680_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	1231 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	199 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/NOT_u1_u1_1435_Update/ca
      -- 
    ca_7345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1435_inst_ack_1, ack => minSumDecode_CP_6680_elements(201)); -- 
    -- CP-element group 202:  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	129 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_exit/$entry
      -- 
    minSumDecode_CP_6680_elements(202) <= minSumDecode_CP_6680_elements(129);
    -- CP-element group 203:  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_exit/$exit
      -- CP-element group 203: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_exit/ack
      -- 
    ack_7349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1381_branch_ack_0, ack => minSumDecode_CP_6680_elements(203)); -- 
    -- CP-element group 204:  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	129 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_taken/$entry
      -- 
    minSumDecode_CP_6680_elements(204) <= minSumDecode_CP_6680_elements(129);
    -- CP-element group 205:  transition  input  no-bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_taken/$exit
      -- CP-element group 205: 	 branch_block_stmt_1353/do_while_stmt_1381/loop_taken/ack
      -- 
    ack_7353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1381_branch_ack_1, ack => minSumDecode_CP_6680_elements(205)); -- 
    -- CP-element group 206:  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	127 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	8 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_1353/do_while_stmt_1381/$exit
      -- 
    minSumDecode_CP_6680_elements(206) <= minSumDecode_CP_6680_elements(127);
    -- CP-element group 207:  transition  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	8 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_1353/if_stmt_1439_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(207) <= minSumDecode_CP_6680_elements(8);
    -- CP-element group 208:  transition  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	8 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_1353/if_stmt_1439_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_1353/if_stmt_1439_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_1353/if_stmt_1439_eval_test/branch_req
      -- 
    branch_req_7362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(208), ack => if_stmt_1439_branch_req_0); -- 
    minSumDecode_CP_6680_elements(208) <= minSumDecode_CP_6680_elements(8);
    -- CP-element group 209:  branch  place  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	212 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_1353/R_bbx_xnphx_xi_readCodeBlockx_xexit_taken_1440_place
      -- 
    minSumDecode_CP_6680_elements(209) <= minSumDecode_CP_6680_elements(208);
    -- CP-element group 210:  transition  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_1353/if_stmt_1439_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(210) <= minSumDecode_CP_6680_elements(209);
    -- CP-element group 211:  transition  input  no-bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	214 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_1353/if_stmt_1439_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_1353/if_stmt_1439_if_link/if_choice_transition
      -- 
    if_choice_transition_7367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1439_branch_ack_1, ack => minSumDecode_CP_6680_elements(211)); -- 
    -- CP-element group 212:  transition  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	209 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_1353/if_stmt_1439_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(212) <= minSumDecode_CP_6680_elements(209);
    -- CP-element group 213:  transition  input  no-bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	9 
    -- CP-element group 213:  members (2) 
      -- CP-element group 213: 	 branch_block_stmt_1353/if_stmt_1439_else_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_1353/if_stmt_1439_else_link/else_choice_transition
      -- 
    else_choice_transition_7371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1439_branch_ack_0, ack => minSumDecode_CP_6680_elements(213)); -- 
    -- CP-element group 214:  place  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	211 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	870 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit
      -- 
    minSumDecode_CP_6680_elements(214) <= minSumDecode_CP_6680_elements(211);
    -- CP-element group 215:  fork  transition  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	10 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (7) 
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/$entry
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_update_start_
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Sample/rr
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Update/cr
      -- 
    rr_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(215), ack => EQ_u16_u1_1453_inst_req_0); -- 
    cr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(215), ack => EQ_u16_u1_1453_inst_req_1); -- 
    minSumDecode_CP_6680_elements(215) <= minSumDecode_CP_6680_elements(10);
    -- CP-element group 216:  transition  input  no-bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Sample/ra
      -- 
    ra_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1453_inst_ack_0, ack => minSumDecode_CP_6680_elements(216)); -- 
    -- CP-element group 217:  transition  input  no-bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	11 
    -- CP-element group 217:  members (4) 
      -- CP-element group 217: 	 branch_block_stmt_1353/assign_stmt_1454/$exit
      -- CP-element group 217: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_1353/assign_stmt_1454/EQ_u16_u1_1453_Update/ca
      -- 
    ca_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1453_inst_ack_1, ack => minSumDecode_CP_6680_elements(217)); -- 
    -- CP-element group 218:  transition  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	11 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 branch_block_stmt_1353/if_stmt_1455_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(218) <= minSumDecode_CP_6680_elements(11);
    -- CP-element group 219:  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	11 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_1353/if_stmt_1455_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_1353/if_stmt_1455_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_1353/if_stmt_1455_eval_test/branch_req
      -- 
    branch_req_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(219), ack => if_stmt_1455_branch_req_0); -- 
    minSumDecode_CP_6680_elements(219) <= minSumDecode_CP_6680_elements(11);
    -- CP-element group 220:  branch  place  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_1353/R_iNsTr_38_1456_place
      -- 
    minSumDecode_CP_6680_elements(220) <= minSumDecode_CP_6680_elements(219);
    -- CP-element group 221:  transition  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_1353/if_stmt_1455_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(221) <= minSumDecode_CP_6680_elements(220);
    -- CP-element group 222:  transition  input  no-bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	225 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_1353/if_stmt_1455_if_link/$exit
      -- CP-element group 222: 	 branch_block_stmt_1353/if_stmt_1455_if_link/if_choice_transition
      -- 
    if_choice_transition_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1455_branch_ack_1, ack => minSumDecode_CP_6680_elements(222)); -- 
    -- CP-element group 223:  transition  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_1353/if_stmt_1455_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(223) <= minSumDecode_CP_6680_elements(220);
    -- CP-element group 224:  transition  input  no-bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_1353/if_stmt_1455_else_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_1353/if_stmt_1455_else_link/else_choice_transition
      -- 
    else_choice_transition_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1455_branch_ack_0, ack => minSumDecode_CP_6680_elements(224)); -- 
    -- CP-element group 225:  place  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	222 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	900 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit
      -- 
    minSumDecode_CP_6680_elements(225) <= minSumDecode_CP_6680_elements(222);
    -- CP-element group 226:  place  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	877 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_1353/readCodeBlockx_xexit_bbx_xnphx_xi1
      -- 
    minSumDecode_CP_6680_elements(226) <= minSumDecode_CP_6680_elements(224);
    -- CP-element group 227:  fork  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	12 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227: 	229 
    -- CP-element group 227: 	230 
    -- CP-element group 227: 	231 
    -- CP-element group 227: 	234 
    -- CP-element group 227: 	235 
    -- CP-element group 227: 	236 
    -- CP-element group 227: 	237 
    -- CP-element group 227: 	238 
    -- CP-element group 227: 	240 
    -- CP-element group 227: 	242 
    -- CP-element group 227: 	245 
    -- CP-element group 227:  members (49) 
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_word_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/word_0/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/word_0/rr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/word_0/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/word_0/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_word_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/word_0/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/word_0/rr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/word_0/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/word_0/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_update_start_
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_complete/$entry
      -- CP-element group 227: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_complete/req
      -- 
    cr_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => LOAD_ebbyNo_1463_load_0_req_1); -- 
    rr_7427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => LOAD_ebbyNo_1463_load_0_req_0); -- 
    cr_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => LOAD_rate_1466_load_0_req_1); -- 
    rr_7460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => LOAD_rate_1466_load_0_req_0); -- 
    cr_7490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => MUL_f32_f32_1471_inst_req_1); -- 
    rr_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => UGT_u16_u1_1477_inst_req_0); -- 
    cr_7504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => UGT_u16_u1_1477_inst_req_1); -- 
    rr_7513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => ADD_u16_u16_1483_inst_req_0); -- 
    cr_7518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => ADD_u16_u16_1483_inst_req_1); -- 
    cr_7532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => type_cast_1487_inst_req_1); -- 
    cr_7546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => ADD_u64_u64_1493_inst_req_1); -- 
    req_7560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(227), ack => MUX_1500_inst_req_1); -- 
    minSumDecode_CP_6680_elements(227) <= minSumDecode_CP_6680_elements(12);
    -- CP-element group 228:  transition  input  no-bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/$exit
      -- CP-element group 228: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Sample/word_access_start/word_0/ra
      -- 
    ra_7428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ebbyNo_1463_load_0_ack_0, ack => minSumDecode_CP_6680_elements(228)); -- 
    -- CP-element group 229:  transition  input  no-bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	232 
    -- CP-element group 229:  members (9) 
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/word_0/$exit
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/word_access_complete/word_0/ca
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/LOAD_ebbyNo_1463_Merge/$entry
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/LOAD_ebbyNo_1463_Merge/$exit
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/LOAD_ebbyNo_1463_Merge/merge_req
      -- CP-element group 229: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_ebbyNo_1463_Update/LOAD_ebbyNo_1463_Merge/merge_ack
      -- 
    ca_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ebbyNo_1463_load_0_ack_1, ack => minSumDecode_CP_6680_elements(229)); -- 
    -- CP-element group 230:  transition  input  no-bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	227 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Sample/word_access_start/word_0/ra
      -- 
    ra_7461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_rate_1466_load_0_ack_0, ack => minSumDecode_CP_6680_elements(230)); -- 
    -- CP-element group 231:  transition  input  no-bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	227 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (9) 
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/word_access_complete/word_0/ca
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/LOAD_rate_1466_Merge/$entry
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/LOAD_rate_1466_Merge/$exit
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/LOAD_rate_1466_Merge/merge_req
      -- CP-element group 231: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/LOAD_rate_1466_Update/LOAD_rate_1466_Merge/merge_ack
      -- 
    ca_7472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_rate_1466_load_0_ack_1, ack => minSumDecode_CP_6680_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	229 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Sample/rr
      -- 
    rr_7485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(232), ack => MUL_f32_f32_1471_inst_req_0); -- 
    minSumDecode_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(229) & minSumDecode_CP_6680_elements(231);
      gj_minSumDecode_cp_element_group_232 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  no-bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Sample/ra
      -- 
    ra_7486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1471_inst_ack_0, ack => minSumDecode_CP_6680_elements(233)); -- 
    -- CP-element group 234:  transition  input  no-bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	227 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	246 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUL_f32_f32_1471_Update/ca
      -- 
    ca_7491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1471_inst_ack_1, ack => minSumDecode_CP_6680_elements(234)); -- 
    -- CP-element group 235:  transition  input  no-bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	227 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Sample/ra
      -- 
    ra_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1477_inst_ack_0, ack => minSumDecode_CP_6680_elements(235)); -- 
    -- CP-element group 236:  transition  input  no-bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	227 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	243 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/UGT_u16_u1_1477_Update/ca
      -- 
    ca_7505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1477_inst_ack_1, ack => minSumDecode_CP_6680_elements(236)); -- 
    -- CP-element group 237:  transition  input  no-bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	227 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Sample/ra
      -- 
    ra_7514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1483_inst_ack_0, ack => minSumDecode_CP_6680_elements(237)); -- 
    -- CP-element group 238:  transition  input  output  no-bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	227 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u16_u16_1483_Update/ca
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Sample/rr
      -- 
    ca_7519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1483_inst_ack_1, ack => minSumDecode_CP_6680_elements(238)); -- 
    rr_7527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(238), ack => type_cast_1487_inst_req_0); -- 
    -- CP-element group 239:  transition  input  no-bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Sample/ra
      -- 
    ra_7528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_0, ack => minSumDecode_CP_6680_elements(239)); -- 
    -- CP-element group 240:  transition  input  output  no-bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	227 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/type_cast_1487_Update/ca
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Sample/rr
      -- 
    ca_7533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_1, ack => minSumDecode_CP_6680_elements(240)); -- 
    rr_7541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(240), ack => ADD_u64_u64_1493_inst_req_0); -- 
    -- CP-element group 241:  transition  input  no-bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Sample/ra
      -- 
    ra_7542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1493_inst_ack_0, ack => minSumDecode_CP_6680_elements(241)); -- 
    -- CP-element group 242:  transition  input  no-bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	227 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/ADD_u64_u64_1493_Update/ca
      -- 
    ca_7547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1493_inst_ack_1, ack => minSumDecode_CP_6680_elements(242)); -- 
    -- CP-element group 243:  join  transition  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	236 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_start/$entry
      -- CP-element group 243: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_start/req
      -- 
    req_7555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(243), ack => MUX_1500_inst_req_0); -- 
    minSumDecode_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(236) & minSumDecode_CP_6680_elements(242);
      gj_minSumDecode_cp_element_group_243 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  transition  input  no-bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_start/$exit
      -- CP-element group 244: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_start/ack
      -- 
    ack_7556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1500_inst_ack_0, ack => minSumDecode_CP_6680_elements(244)); -- 
    -- CP-element group 245:  transition  input  no-bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	227 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_complete/$exit
      -- CP-element group 245: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/MUX_1500_complete/ack
      -- 
    ack_7561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1500_inst_ack_1, ack => minSumDecode_CP_6680_elements(245)); -- 
    -- CP-element group 246:  join  transition  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	234 
    -- CP-element group 246: 	244 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	13 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_1353/assign_stmt_1464_to_assign_stmt_1501/$exit
      -- 
    minSumDecode_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(234) & minSumDecode_CP_6680_elements(244) & minSumDecode_CP_6680_elements(245);
      gj_minSumDecode_cp_element_group_246 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	14 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247: 	249 
    -- CP-element group 247: 	250 
    -- CP-element group 247: 	251 
    -- CP-element group 247: 	253 
    -- CP-element group 247: 	255 
    -- CP-element group 247: 	257 
    -- CP-element group 247: 	260 
    -- CP-element group 247: 	261 
    -- CP-element group 247: 	262 
    -- CP-element group 247: 	264 
    -- CP-element group 247:  members (80) 
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_scale_0/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_final_index_sum_regn/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_final_index_sum_regn/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_scale_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_resize_0/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_request/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_scale_0/scale_rename_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_final_index_sum_regn/ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_base_plus_offset/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_complete/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_base_plus_offset/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_base_plus_offset/sum_rename_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_final_index_sum_regn/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_scale_0/scale_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_base_plus_offset/sum_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_request/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_resize_0/index_resize_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_resize_0/index_resize_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_root_address_calculated
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_offset_calculated
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_resized_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_scaled_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_computed_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_resize_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_resize_0/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_resize_0/index_resize_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_resize_0/index_resize_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_scale_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_scale_0/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_scale_0/scale_rename_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_index_scale_0/scale_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_final_index_sum_regn/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_final_index_sum_regn/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_final_index_sum_regn/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_final_index_sum_regn/ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_base_plus_offset/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_base_plus_offset/$exit
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_base_plus_offset/sum_rename_req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1514_base_plus_offset/sum_rename_ack
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_request/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_request/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_complete/req
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_root_address_calculated
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_offset_calculated
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_resized_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_scaled_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_computed_0
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/array_obj_ref_1519_index_resize_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/word_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/word_0/cr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/word_0/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/word_0/cr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Sample/rr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Update/cr
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Update/cr
      -- 
    req_7602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => addr_of_1515_final_reg_req_1); -- 
    req_7597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => addr_of_1515_final_reg_req_0); -- 
    req_7641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => addr_of_1520_final_reg_req_1); -- 
    req_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => addr_of_1520_final_reg_req_0); -- 
    cr_7686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => ptr_deref_1524_load_0_req_1); -- 
    cr_7705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => MUL_f32_f32_1530_inst_req_1); -- 
    cr_7719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => MUL_f32_f32_1535_inst_req_1); -- 
    cr_7769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => ptr_deref_1538_store_0_req_1); -- 
    rr_7778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => ADD_u64_u64_1545_inst_req_0); -- 
    cr_7783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => ADD_u64_u64_1545_inst_req_1); -- 
    cr_7797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(247), ack => EQ_u64_u1_1550_inst_req_1); -- 
    minSumDecode_CP_6680_elements(247) <= minSumDecode_CP_6680_elements(14);
    -- CP-element group 248:  transition  input  no-bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	265 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_request/$exit
      -- CP-element group 248: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_request/ack
      -- 
    ack_7598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1515_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (24) 
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_complete/$exit
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1515_complete/ack
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_word_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_address_resized
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_addr_resize/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_addr_resize/$exit
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_addr_resize/base_resize_req
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_addr_resize/base_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_word_addrgen/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_word_addrgen/$exit
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_word_addrgen/root_register_req
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_word_addrgen/root_register_ack
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/word_0/rr
      -- 
    ack_7603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1515_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(249)); -- 
    rr_7675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(249), ack => ptr_deref_1524_load_0_req_0); -- 
    -- CP-element group 250:  transition  input  no-bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	247 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	265 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_request/$exit
      -- CP-element group 250: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_request/ack
      -- CP-element group 250: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_sample_completed_
      -- 
    ack_7637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1520_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  no-bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	247 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	258 
    -- CP-element group 251:  members (19) 
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_complete/ack
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_complete/$exit
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/addr_of_1520_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_word_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_root_address_calculated
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_address_resized
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_addr_resize/$entry
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_addr_resize/$exit
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_addr_resize/base_resize_req
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_addr_resize/base_resize_ack
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_plus_offset/$entry
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_plus_offset/$exit
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_plus_offset/sum_rename_req
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_base_plus_offset/sum_rename_ack
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_word_addrgen/$entry
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_word_addrgen/$exit
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_word_addrgen/root_register_req
      -- CP-element group 251: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_word_addrgen/root_register_ack
      -- 
    ack_7642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1520_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(251)); -- 
    -- CP-element group 252:  transition  input  no-bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (5) 
      -- CP-element group 252: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/$exit
      -- CP-element group 252: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/word_0/$exit
      -- CP-element group 252: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Sample/word_access_start/word_0/ra
      -- 
    ra_7676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1524_load_0_ack_0, ack => minSumDecode_CP_6680_elements(252)); -- 
    -- CP-element group 253:  transition  input  output  no-bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	247 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (12) 
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/$exit
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/word_0/$exit
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/word_access_complete/word_0/ca
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/ptr_deref_1524_Merge/$entry
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/ptr_deref_1524_Merge/$exit
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/ptr_deref_1524_Merge/merge_req
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1524_Update/ptr_deref_1524_Merge/merge_ack
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Sample/rr
      -- 
    ca_7687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1524_load_0_ack_1, ack => minSumDecode_CP_6680_elements(253)); -- 
    rr_7700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(253), ack => MUL_f32_f32_1530_inst_req_0); -- 
    -- CP-element group 254:  transition  input  no-bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Sample/ra
      -- 
    ra_7701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1530_inst_ack_0, ack => minSumDecode_CP_6680_elements(254)); -- 
    -- CP-element group 255:  transition  input  output  no-bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	247 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1530_Update/ca
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Sample/rr
      -- 
    ca_7706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1530_inst_ack_1, ack => minSumDecode_CP_6680_elements(255)); -- 
    rr_7714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(255), ack => MUL_f32_f32_1535_inst_req_0); -- 
    -- CP-element group 256:  transition  input  no-bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Sample/ra
      -- 
    ra_7715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1535_inst_ack_0, ack => minSumDecode_CP_6680_elements(256)); -- 
    -- CP-element group 257:  transition  input  no-bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	247 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/MUL_f32_f32_1535_Update/ca
      -- 
    ca_7720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_f32_f32_1535_inst_ack_1, ack => minSumDecode_CP_6680_elements(257)); -- 
    -- CP-element group 258:  join  transition  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	251 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (9) 
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/ptr_deref_1538_Split/$entry
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/ptr_deref_1538_Split/$exit
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/ptr_deref_1538_Split/split_req
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/ptr_deref_1538_Split/split_ack
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/$entry
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/word_0/$entry
      -- CP-element group 258: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/word_0/rr
      -- 
    rr_7758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(258), ack => ptr_deref_1538_store_0_req_0); -- 
    minSumDecode_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(251) & minSumDecode_CP_6680_elements(257);
      gj_minSumDecode_cp_element_group_258 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  transition  input  no-bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (5) 
      -- CP-element group 259: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/$exit
      -- CP-element group 259: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/word_0/$exit
      -- CP-element group 259: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Sample/word_access_start/word_0/ra
      -- 
    ra_7759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1538_store_0_ack_0, ack => minSumDecode_CP_6680_elements(259)); -- 
    -- CP-element group 260:  transition  input  no-bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	247 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	265 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/$exit
      -- CP-element group 260: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/word_0/$exit
      -- CP-element group 260: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ptr_deref_1538_Update/word_access_complete/word_0/ca
      -- 
    ca_7770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1538_store_0_ack_1, ack => minSumDecode_CP_6680_elements(260)); -- 
    -- CP-element group 261:  transition  input  no-bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	247 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Sample/ra
      -- 
    ra_7779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1545_inst_ack_0, ack => minSumDecode_CP_6680_elements(261)); -- 
    -- CP-element group 262:  transition  input  output  no-bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	247 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/ADD_u64_u64_1545_Update/ca
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Sample/rr
      -- 
    ca_7784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1545_inst_ack_1, ack => minSumDecode_CP_6680_elements(262)); -- 
    rr_7792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(262), ack => EQ_u64_u1_1550_inst_req_0); -- 
    -- CP-element group 263:  transition  input  no-bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Sample/ra
      -- 
    ra_7793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1550_inst_ack_0, ack => minSumDecode_CP_6680_elements(263)); -- 
    -- CP-element group 264:  transition  input  no-bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	247 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/EQ_u64_u1_1550_Update/ca
      -- 
    ca_7798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1550_inst_ack_1, ack => minSumDecode_CP_6680_elements(264)); -- 
    -- CP-element group 265:  join  transition  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	248 
    -- CP-element group 265: 	250 
    -- CP-element group 265: 	260 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	15 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_1353/assign_stmt_1516_to_assign_stmt_1551/$exit
      -- 
    minSumDecode_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(248) & minSumDecode_CP_6680_elements(250) & minSumDecode_CP_6680_elements(260) & minSumDecode_CP_6680_elements(264);
      gj_minSumDecode_cp_element_group_265 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	15 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (1) 
      -- CP-element group 266: 	 branch_block_stmt_1353/if_stmt_1552_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(266) <= minSumDecode_CP_6680_elements(15);
    -- CP-element group 267:  transition  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	15 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1353/if_stmt_1552_eval_test/$entry
      -- CP-element group 267: 	 branch_block_stmt_1353/if_stmt_1552_eval_test/$exit
      -- CP-element group 267: 	 branch_block_stmt_1353/if_stmt_1552_eval_test/branch_req
      -- 
    branch_req_7806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(267), ack => if_stmt_1552_branch_req_0); -- 
    minSumDecode_CP_6680_elements(267) <= minSumDecode_CP_6680_elements(15);
    -- CP-element group 268:  branch  place  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	271 
    -- CP-element group 268:  members (1) 
      -- CP-element group 268: 	 branch_block_stmt_1353/R_exitcond_1553_place
      -- 
    minSumDecode_CP_6680_elements(268) <= minSumDecode_CP_6680_elements(267);
    -- CP-element group 269:  transition  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (1) 
      -- CP-element group 269: 	 branch_block_stmt_1353/if_stmt_1552_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(269) <= minSumDecode_CP_6680_elements(268);
    -- CP-element group 270:  transition  input  no-bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	273 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_1353/if_stmt_1552_if_link/$exit
      -- CP-element group 270: 	 branch_block_stmt_1353/if_stmt_1552_if_link/if_choice_transition
      -- 
    if_choice_transition_7811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1552_branch_ack_1, ack => minSumDecode_CP_6680_elements(270)); -- 
    -- CP-element group 271:  transition  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (1) 
      -- CP-element group 271: 	 branch_block_stmt_1353/if_stmt_1552_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(271) <= minSumDecode_CP_6680_elements(268);
    -- CP-element group 272:  transition  input  no-bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (2) 
      -- CP-element group 272: 	 branch_block_stmt_1353/if_stmt_1552_else_link/$exit
      -- CP-element group 272: 	 branch_block_stmt_1353/if_stmt_1552_else_link/else_choice_transition
      -- 
    else_choice_transition_7815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1552_branch_ack_0, ack => minSumDecode_CP_6680_elements(272)); -- 
    -- CP-element group 273:  place  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	270 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	890 
    -- CP-element group 273:  members (1) 
      -- CP-element group 273: 	 branch_block_stmt_1353/bb_6_initialize_aPriorix_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(273) <= minSumDecode_CP_6680_elements(270);
    -- CP-element group 274:  place  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	880 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_1353/bb_6_bb_6
      -- 
    minSumDecode_CP_6680_elements(274) <= minSumDecode_CP_6680_elements(272);
    -- CP-element group 275:  fork  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	17 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: 	277 
    -- CP-element group 275: 	279 
    -- CP-element group 275:  members (16) 
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_update_start_
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_word_address_calculated
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_root_address_calculated
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/word_0/rr
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/word_0/cr
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_update_start_
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Update/cr
      -- 
    cr_7847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(275), ack => LOAD_ncol_ind_1573_load_0_req_1); -- 
    rr_7836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(275), ack => LOAD_ncol_ind_1573_load_0_req_0); -- 
    cr_7866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(275), ack => EQ_u16_u1_1579_inst_req_1); -- 
    minSumDecode_CP_6680_elements(275) <= minSumDecode_CP_6680_elements(17);
    -- CP-element group 276:  transition  input  no-bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/$exit
      -- CP-element group 276: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/word_0/$exit
      -- CP-element group 276: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Sample/word_access_start/word_0/ra
      -- 
    ra_7837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_1573_load_0_ack_0, ack => minSumDecode_CP_6680_elements(276)); -- 
    -- CP-element group 277:  transition  input  output  no-bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (12) 
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/$exit
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/word_0/$exit
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/word_access_complete/word_0/ca
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/LOAD_ncol_ind_1573_Merge/$entry
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/LOAD_ncol_ind_1573_Merge/$exit
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/LOAD_ncol_ind_1573_Merge/merge_req
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/LOAD_ncol_ind_1573_Update/LOAD_ncol_ind_1573_Merge/merge_ack
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Sample/rr
      -- 
    ca_7848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_1573_load_0_ack_1, ack => minSumDecode_CP_6680_elements(277)); -- 
    rr_7861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(277), ack => EQ_u16_u1_1579_inst_req_0); -- 
    -- CP-element group 278:  transition  input  no-bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Sample/ra
      -- 
    ra_7862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1579_inst_ack_0, ack => minSumDecode_CP_6680_elements(278)); -- 
    -- CP-element group 279:  transition  input  no-bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	275 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	18 
    -- CP-element group 279:  members (4) 
      -- CP-element group 279: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/$exit
      -- CP-element group 279: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_1353/assign_stmt_1574_to_assign_stmt_1580/EQ_u16_u1_1579_Update/ca
      -- 
    ca_7867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1579_inst_ack_1, ack => minSumDecode_CP_6680_elements(279)); -- 
    -- CP-element group 280:  transition  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	18 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_1353/if_stmt_1581_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(280) <= minSumDecode_CP_6680_elements(18);
    -- CP-element group 281:  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	18 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1353/if_stmt_1581_eval_test/$entry
      -- CP-element group 281: 	 branch_block_stmt_1353/if_stmt_1581_eval_test/$exit
      -- CP-element group 281: 	 branch_block_stmt_1353/if_stmt_1581_eval_test/branch_req
      -- 
    branch_req_7875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(281), ack => if_stmt_1581_branch_req_0); -- 
    minSumDecode_CP_6680_elements(281) <= minSumDecode_CP_6680_elements(18);
    -- CP-element group 282:  branch  place  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: 	285 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_1353/R_iNsTr_7_1582_place
      -- 
    minSumDecode_CP_6680_elements(282) <= minSumDecode_CP_6680_elements(281);
    -- CP-element group 283:  transition  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_1353/if_stmt_1581_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(283) <= minSumDecode_CP_6680_elements(282);
    -- CP-element group 284:  transition  input  no-bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	287 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_1353/if_stmt_1581_if_link/$exit
      -- CP-element group 284: 	 branch_block_stmt_1353/if_stmt_1581_if_link/if_choice_transition
      -- 
    if_choice_transition_7880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1581_branch_ack_1, ack => minSumDecode_CP_6680_elements(284)); -- 
    -- CP-element group 285:  transition  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	282 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_1353/if_stmt_1581_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(285) <= minSumDecode_CP_6680_elements(282);
    -- CP-element group 286:  transition  input  no-bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_1353/if_stmt_1581_else_link/$exit
      -- CP-element group 286: 	 branch_block_stmt_1353/if_stmt_1581_else_link/else_choice_transition
      -- 
    else_choice_transition_7884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1581_branch_ack_0, ack => minSumDecode_CP_6680_elements(286)); -- 
    -- CP-element group 287:  place  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	284 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	926 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader
      -- 
    minSumDecode_CP_6680_elements(287) <= minSumDecode_CP_6680_elements(284);
    -- CP-element group 288:  place  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	906 
    -- CP-element group 288:  members (1) 
      -- CP-element group 288: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_bbx_xnphx_xi5
      -- 
    minSumDecode_CP_6680_elements(288) <= minSumDecode_CP_6680_elements(286);
    -- CP-element group 289:  fork  transition  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	19 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289: 	291 
    -- CP-element group 289: 	292 
    -- CP-element group 289: 	293 
    -- CP-element group 289: 	295 
    -- CP-element group 289: 	297 
    -- CP-element group 289: 	300 
    -- CP-element group 289:  members (22) 
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_update_start_
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_complete/$entry
      -- CP-element group 289: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_complete/req
      -- 
    rr_7897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => UGT_u16_u1_1592_inst_req_0); -- 
    cr_7902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => UGT_u16_u1_1592_inst_req_1); -- 
    rr_7911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => ADD_u16_u16_1598_inst_req_0); -- 
    cr_7916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => ADD_u16_u16_1598_inst_req_1); -- 
    cr_7930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => type_cast_1602_inst_req_1); -- 
    cr_7944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => ADD_u64_u64_1608_inst_req_1); -- 
    req_7958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(289), ack => MUX_1615_inst_req_1); -- 
    minSumDecode_CP_6680_elements(289) <= minSumDecode_CP_6680_elements(19);
    -- CP-element group 290:  transition  input  no-bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Sample/ra
      -- 
    ra_7898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1592_inst_ack_0, ack => minSumDecode_CP_6680_elements(290)); -- 
    -- CP-element group 291:  transition  input  no-bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	298 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/UGT_u16_u1_1592_Update/ca
      -- 
    ca_7903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1592_inst_ack_1, ack => minSumDecode_CP_6680_elements(291)); -- 
    -- CP-element group 292:  transition  input  no-bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	289 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Sample/ra
      -- 
    ra_7912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1598_inst_ack_0, ack => minSumDecode_CP_6680_elements(292)); -- 
    -- CP-element group 293:  transition  input  output  no-bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	289 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u16_u16_1598_Update/ca
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Sample/rr
      -- 
    ca_7917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1598_inst_ack_1, ack => minSumDecode_CP_6680_elements(293)); -- 
    rr_7925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(293), ack => type_cast_1602_inst_req_0); -- 
    -- CP-element group 294:  transition  input  no-bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Sample/ra
      -- 
    ra_7926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1602_inst_ack_0, ack => minSumDecode_CP_6680_elements(294)); -- 
    -- CP-element group 295:  transition  input  output  no-bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	289 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/type_cast_1602_Update/ca
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Sample/rr
      -- 
    ca_7931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1602_inst_ack_1, ack => minSumDecode_CP_6680_elements(295)); -- 
    rr_7939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(295), ack => ADD_u64_u64_1608_inst_req_0); -- 
    -- CP-element group 296:  transition  input  no-bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Sample/ra
      -- 
    ra_7940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1608_inst_ack_0, ack => minSumDecode_CP_6680_elements(296)); -- 
    -- CP-element group 297:  transition  input  no-bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	289 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/ADD_u64_u64_1608_Update/ca
      -- 
    ca_7945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1608_inst_ack_1, ack => minSumDecode_CP_6680_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	291 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_start/$entry
      -- CP-element group 298: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_start/req
      -- 
    req_7953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(298), ack => MUX_1615_inst_req_0); -- 
    minSumDecode_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(291) & minSumDecode_CP_6680_elements(297);
      gj_minSumDecode_cp_element_group_298 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  transition  input  no-bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_start/$exit
      -- CP-element group 299: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_start/ack
      -- 
    ack_7954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1615_inst_ack_0, ack => minSumDecode_CP_6680_elements(299)); -- 
    -- CP-element group 300:  transition  input  no-bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	289 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_complete/$exit
      -- CP-element group 300: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/MUX_1615_complete/ack
      -- 
    ack_7959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1615_inst_ack_1, ack => minSumDecode_CP_6680_elements(300)); -- 
    -- CP-element group 301:  join  transition  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	20 
    -- CP-element group 301:  members (1) 
      -- CP-element group 301: 	 branch_block_stmt_1353/assign_stmt_1593_to_assign_stmt_1616/$exit
      -- 
    minSumDecode_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(299) & minSumDecode_CP_6680_elements(300);
      gj_minSumDecode_cp_element_group_301 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	21 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302: 	304 
    -- CP-element group 302: 	305 
    -- CP-element group 302: 	306 
    -- CP-element group 302: 	308 
    -- CP-element group 302: 	310 
    -- CP-element group 302: 	312 
    -- CP-element group 302: 	314 
    -- CP-element group 302: 	316 
    -- CP-element group 302: 	318 
    -- CP-element group 302: 	321 
    -- CP-element group 302: 	322 
    -- CP-element group 302: 	323 
    -- CP-element group 302: 	325 
    -- CP-element group 302:  members (70) 
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_root_address_calculated
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_offset_calculated
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_resized_0
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_scaled_0
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_computed_0
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_resize_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_resize_0/$exit
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_resize_0/index_resize_req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_resize_0/index_resize_ack
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_scale_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_scale_0/$exit
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_scale_0/scale_rename_req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_index_scale_0/scale_rename_ack
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_final_index_sum_regn/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_final_index_sum_regn/$exit
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_final_index_sum_regn/req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_final_index_sum_regn/ack
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_base_plus_offset/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_base_plus_offset/$exit
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_base_plus_offset/sum_rename_req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1629_base_plus_offset/sum_rename_ack
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_request/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_request/req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_complete/req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_complete/req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/word_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/word_0/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_complete/req
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/word_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/word_0/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/word_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/word_0/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Update/cr
      -- 
    req_8000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => addr_of_1630_final_reg_req_1); -- 
    req_7995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => addr_of_1630_final_reg_req_0); -- 
    rr_8009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ADD_u64_u64_1636_inst_req_0); -- 
    cr_8014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ADD_u64_u64_1636_inst_req_1); -- 
    req_8053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => addr_of_1641_final_reg_req_1); -- 
    cr_8098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ptr_deref_1645_load_0_req_1); -- 
    cr_8117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ADD_u16_u16_1651_inst_req_1); -- 
    cr_8131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => type_cast_1655_inst_req_1); -- 
    req_8170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => addr_of_1660_final_reg_req_1); -- 
    cr_8215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ptr_deref_1664_load_0_req_1); -- 
    cr_8270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ptr_deref_1667_store_0_req_1); -- 
    rr_8279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ADD_u64_u64_1674_inst_req_0); -- 
    cr_8284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => ADD_u64_u64_1674_inst_req_1); -- 
    cr_8298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(302), ack => EQ_u64_u1_1679_inst_req_1); -- 
    minSumDecode_CP_6680_elements(302) <= minSumDecode_CP_6680_elements(21);
    -- CP-element group 303:  transition  input  no-bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	326 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_request/$exit
      -- CP-element group 303: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_request/ack
      -- 
    ack_7996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1630_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  no-bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	319 
    -- CP-element group 304:  members (19) 
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_complete/$exit
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1630_complete/ack
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_address_calculated
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_word_address_calculated
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_root_address_calculated
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_address_resized
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_addr_resize/$entry
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_addr_resize/$exit
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_addr_resize/base_resize_req
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_addr_resize/base_resize_ack
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_plus_offset/$entry
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_plus_offset/$exit
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_plus_offset/sum_rename_req
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_base_plus_offset/sum_rename_ack
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_word_addrgen/$entry
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_word_addrgen/$exit
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_word_addrgen/root_register_req
      -- CP-element group 304: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_word_addrgen/root_register_ack
      -- 
    ack_8001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1630_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(304)); -- 
    -- CP-element group 305:  transition  input  no-bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	302 
    -- CP-element group 305: successors 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Sample/ra
      -- 
    ra_8010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1636_inst_ack_0, ack => minSumDecode_CP_6680_elements(305)); -- 
    -- CP-element group 306:  transition  input  output  no-bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	302 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (27) 
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1636_Update/ca
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_root_address_calculated
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_offset_calculated
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_resized_0
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_scaled_0
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_computed_0
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_resize_0/$entry
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_resize_0/$exit
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_resize_0/index_resize_req
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_resize_0/index_resize_ack
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_scale_0/$entry
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_scale_0/$exit
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_scale_0/scale_rename_req
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_index_scale_0/scale_rename_ack
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_final_index_sum_regn/$entry
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_final_index_sum_regn/$exit
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_final_index_sum_regn/req
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_final_index_sum_regn/ack
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_base_plus_offset/$entry
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_base_plus_offset/$exit
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_base_plus_offset/sum_rename_req
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1640_base_plus_offset/sum_rename_ack
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_request/$entry
      -- CP-element group 306: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_request/req
      -- 
    ca_8015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1636_inst_ack_1, ack => minSumDecode_CP_6680_elements(306)); -- 
    req_8048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(306), ack => addr_of_1641_final_reg_req_0); -- 
    -- CP-element group 307:  transition  input  no-bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	326 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_request/$exit
      -- CP-element group 307: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_request/ack
      -- 
    ack_8049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1641_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(307)); -- 
    -- CP-element group 308:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	302 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (24) 
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_complete/$exit
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1641_complete/ack
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_address_resized
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_addr_resize/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_addr_resize/$exit
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_addr_resize/base_resize_req
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_addr_resize/base_resize_ack
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_plus_offset/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_plus_offset/$exit
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_plus_offset/sum_rename_req
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_base_plus_offset/sum_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_word_addrgen/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_word_addrgen/$exit
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_word_addrgen/root_register_req
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_word_addrgen/root_register_ack
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/word_0/rr
      -- 
    ack_8054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1641_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(308)); -- 
    rr_8087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(308), ack => ptr_deref_1645_load_0_req_0); -- 
    -- CP-element group 309:  transition  input  no-bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (5) 
      -- CP-element group 309: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/$exit
      -- CP-element group 309: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/word_0/$exit
      -- CP-element group 309: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Sample/word_access_start/word_0/ra
      -- 
    ra_8088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1645_load_0_ack_0, ack => minSumDecode_CP_6680_elements(309)); -- 
    -- CP-element group 310:  transition  input  output  no-bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	302 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (12) 
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/$exit
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/word_0/$exit
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/word_access_complete/word_0/ca
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/ptr_deref_1645_Merge/$entry
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/ptr_deref_1645_Merge/$exit
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/ptr_deref_1645_Merge/merge_req
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1645_Update/ptr_deref_1645_Merge/merge_ack
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Sample/rr
      -- 
    ca_8099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1645_load_0_ack_1, ack => minSumDecode_CP_6680_elements(310)); -- 
    rr_8112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(310), ack => ADD_u16_u16_1651_inst_req_0); -- 
    -- CP-element group 311:  transition  input  no-bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Sample/ra
      -- 
    ra_8113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1651_inst_ack_0, ack => minSumDecode_CP_6680_elements(311)); -- 
    -- CP-element group 312:  transition  input  output  no-bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	302 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u16_u16_1651_Update/ca
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Sample/rr
      -- 
    ca_8118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1651_inst_ack_1, ack => minSumDecode_CP_6680_elements(312)); -- 
    rr_8126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(312), ack => type_cast_1655_inst_req_0); -- 
    -- CP-element group 313:  transition  input  no-bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Sample/ra
      -- 
    ra_8127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1655_inst_ack_0, ack => minSumDecode_CP_6680_elements(313)); -- 
    -- CP-element group 314:  transition  input  output  no-bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	302 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (27) 
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_root_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/type_cast_1655_Update/ca
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_offset_calculated
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_resized_0
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_scaled_0
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_computed_0
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_resize_0/$entry
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_resize_0/$exit
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_resize_0/index_resize_req
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_resize_0/index_resize_ack
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_scale_0/$entry
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_scale_0/$exit
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_scale_0/scale_rename_req
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_index_scale_0/scale_rename_ack
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_final_index_sum_regn/$entry
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_final_index_sum_regn/$exit
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_final_index_sum_regn/req
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_final_index_sum_regn/ack
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_base_plus_offset/$entry
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_base_plus_offset/$exit
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_base_plus_offset/sum_rename_req
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/array_obj_ref_1659_base_plus_offset/sum_rename_ack
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_request/$entry
      -- CP-element group 314: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_request/req
      -- 
    ca_8132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1655_inst_ack_1, ack => minSumDecode_CP_6680_elements(314)); -- 
    req_8165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(314), ack => addr_of_1660_final_reg_req_0); -- 
    -- CP-element group 315:  transition  input  no-bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	326 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_request/$exit
      -- CP-element group 315: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_request/ack
      -- 
    ack_8166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1660_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(315)); -- 
    -- CP-element group 316:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	302 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (24) 
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_complete/$exit
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/addr_of_1660_complete/ack
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_word_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_root_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_address_resized
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_addr_resize/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_addr_resize/$exit
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_addr_resize/base_resize_req
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_addr_resize/base_resize_ack
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_plus_offset/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_plus_offset/$exit
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_plus_offset/sum_rename_req
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_base_plus_offset/sum_rename_ack
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_word_addrgen/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_word_addrgen/$exit
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_word_addrgen/root_register_req
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_word_addrgen/root_register_ack
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/word_0/$entry
      -- CP-element group 316: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/word_0/rr
      -- 
    ack_8171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1660_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(316)); -- 
    rr_8204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(316), ack => ptr_deref_1664_load_0_req_0); -- 
    -- CP-element group 317:  transition  input  no-bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317:  members (5) 
      -- CP-element group 317: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/$exit
      -- CP-element group 317: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/word_0/$exit
      -- CP-element group 317: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Sample/word_access_start/word_0/ra
      -- 
    ra_8205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_load_0_ack_0, ack => minSumDecode_CP_6680_elements(317)); -- 
    -- CP-element group 318:  transition  input  no-bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	302 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (9) 
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/$exit
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/word_0/$exit
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/word_access_complete/word_0/ca
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/ptr_deref_1664_Merge/$entry
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/ptr_deref_1664_Merge/$exit
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/ptr_deref_1664_Merge/merge_req
      -- CP-element group 318: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1664_Update/ptr_deref_1664_Merge/merge_ack
      -- 
    ca_8216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_load_0_ack_1, ack => minSumDecode_CP_6680_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	304 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (9) 
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/ptr_deref_1667_Split/$entry
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/ptr_deref_1667_Split/$exit
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/ptr_deref_1667_Split/split_req
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/ptr_deref_1667_Split/split_ack
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/$entry
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/word_0/$entry
      -- CP-element group 319: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/word_0/rr
      -- 
    rr_8259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(319), ack => ptr_deref_1667_store_0_req_0); -- 
    minSumDecode_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(304) & minSumDecode_CP_6680_elements(318);
      gj_minSumDecode_cp_element_group_319 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  transition  input  no-bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/$exit
      -- CP-element group 320: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/word_0/$exit
      -- CP-element group 320: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Sample/word_access_start/word_0/ra
      -- 
    ra_8260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1667_store_0_ack_0, ack => minSumDecode_CP_6680_elements(320)); -- 
    -- CP-element group 321:  transition  input  no-bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	302 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	326 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/$exit
      -- CP-element group 321: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/word_0/$exit
      -- CP-element group 321: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ptr_deref_1667_Update/word_access_complete/word_0/ca
      -- 
    ca_8271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1667_store_0_ack_1, ack => minSumDecode_CP_6680_elements(321)); -- 
    -- CP-element group 322:  transition  input  no-bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	302 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Sample/ra
      -- 
    ra_8280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1674_inst_ack_0, ack => minSumDecode_CP_6680_elements(322)); -- 
    -- CP-element group 323:  transition  input  output  no-bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	302 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/ADD_u64_u64_1674_Update/ca
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Sample/rr
      -- 
    ca_8285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1674_inst_ack_1, ack => minSumDecode_CP_6680_elements(323)); -- 
    rr_8293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(323), ack => EQ_u64_u1_1679_inst_req_0); -- 
    -- CP-element group 324:  transition  input  no-bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Sample/ra
      -- 
    ra_8294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1679_inst_ack_0, ack => minSumDecode_CP_6680_elements(324)); -- 
    -- CP-element group 325:  transition  input  no-bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	302 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/EQ_u64_u1_1679_Update/ca
      -- 
    ca_8299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1679_inst_ack_1, ack => minSumDecode_CP_6680_elements(325)); -- 
    -- CP-element group 326:  join  transition  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	303 
    -- CP-element group 326: 	307 
    -- CP-element group 326: 	315 
    -- CP-element group 326: 	321 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	22 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_1353/assign_stmt_1631_to_assign_stmt_1680/$exit
      -- 
    minSumDecode_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(303) & minSumDecode_CP_6680_elements(307) & minSumDecode_CP_6680_elements(315) & minSumDecode_CP_6680_elements(321) & minSumDecode_CP_6680_elements(325);
      gj_minSumDecode_cp_element_group_326 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	22 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (1) 
      -- CP-element group 327: 	 branch_block_stmt_1353/if_stmt_1681_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(327) <= minSumDecode_CP_6680_elements(22);
    -- CP-element group 328:  transition  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	22 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_1353/if_stmt_1681_eval_test/$entry
      -- CP-element group 328: 	 branch_block_stmt_1353/if_stmt_1681_eval_test/$exit
      -- CP-element group 328: 	 branch_block_stmt_1353/if_stmt_1681_eval_test/branch_req
      -- 
    branch_req_8307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(328), ack => if_stmt_1681_branch_req_0); -- 
    minSumDecode_CP_6680_elements(328) <= minSumDecode_CP_6680_elements(22);
    -- CP-element group 329:  branch  place  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329: 	332 
    -- CP-element group 329:  members (1) 
      -- CP-element group 329: 	 branch_block_stmt_1353/R_exitcond3_1682_place
      -- 
    minSumDecode_CP_6680_elements(329) <= minSumDecode_CP_6680_elements(328);
    -- CP-element group 330:  transition  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_1353/if_stmt_1681_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(330) <= minSumDecode_CP_6680_elements(329);
    -- CP-element group 331:  transition  input  no-bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	334 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_1353/if_stmt_1681_if_link/$exit
      -- CP-element group 331: 	 branch_block_stmt_1353/if_stmt_1681_if_link/if_choice_transition
      -- 
    if_choice_transition_8312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1681_branch_ack_1, ack => minSumDecode_CP_6680_elements(331)); -- 
    -- CP-element group 332:  transition  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	329 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (1) 
      -- CP-element group 332: 	 branch_block_stmt_1353/if_stmt_1681_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(332) <= minSumDecode_CP_6680_elements(329);
    -- CP-element group 333:  transition  input  no-bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_1353/if_stmt_1681_else_link/$exit
      -- CP-element group 333: 	 branch_block_stmt_1353/if_stmt_1681_else_link/else_choice_transition
      -- 
    else_choice_transition_8316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1681_branch_ack_0, ack => minSumDecode_CP_6680_elements(333)); -- 
    -- CP-element group 334:  place  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	331 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	919 
    -- CP-element group 334:  members (1) 
      -- CP-element group 334: 	 branch_block_stmt_1353/bb_10_initializeMessagex_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(334) <= minSumDecode_CP_6680_elements(331);
    -- CP-element group 335:  place  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	909 
    -- CP-element group 335:  members (1) 
      -- CP-element group 335: 	 branch_block_stmt_1353/bb_10_bb_10
      -- 
    minSumDecode_CP_6680_elements(335) <= minSumDecode_CP_6680_elements(333);
    -- CP-element group 336:  fork  transition  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	25 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	338 
    -- CP-element group 336: 	339 
    -- CP-element group 336: 	340 
    -- CP-element group 336: 	343 
    -- CP-element group 336:  members (22) 
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_update_start_
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Sample/rr
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Update/cr
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_update_start_
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_word_address_calculated
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_root_address_calculated
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/word_0/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/word_0/rr
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/word_0/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/word_0/cr
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_update_start_
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Update/cr
      -- 
    rr_8329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(336), ack => ADD_u16_u16_1724_inst_req_0); -- 
    cr_8334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(336), ack => ADD_u16_u16_1724_inst_req_1); -- 
    cr_8362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(336), ack => LOAD_maxNitr_1727_load_0_req_1); -- 
    rr_8351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(336), ack => LOAD_maxNitr_1727_load_0_req_0); -- 
    cr_8381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(336), ack => ULT_u16_u1_1732_inst_req_1); -- 
    minSumDecode_CP_6680_elements(336) <= minSumDecode_CP_6680_elements(25);
    -- CP-element group 337:  transition  input  no-bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Sample/ra
      -- 
    ra_8330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1724_inst_ack_0, ack => minSumDecode_CP_6680_elements(337)); -- 
    -- CP-element group 338:  transition  input  no-bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	341 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ADD_u16_u16_1724_Update/ca
      -- 
    ca_8335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1724_inst_ack_1, ack => minSumDecode_CP_6680_elements(338)); -- 
    -- CP-element group 339:  transition  input  no-bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	336 
    -- CP-element group 339: successors 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/$exit
      -- CP-element group 339: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/word_0/$exit
      -- CP-element group 339: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Sample/word_access_start/word_0/ra
      -- 
    ra_8352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_maxNitr_1727_load_0_ack_0, ack => minSumDecode_CP_6680_elements(339)); -- 
    -- CP-element group 340:  transition  input  no-bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	336 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (9) 
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/$exit
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/word_access_complete/word_0/ca
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/LOAD_maxNitr_1727_Merge/$entry
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/LOAD_maxNitr_1727_Merge/$exit
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/LOAD_maxNitr_1727_Merge/merge_req
      -- CP-element group 340: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/LOAD_maxNitr_1727_Update/LOAD_maxNitr_1727_Merge/merge_ack
      -- 
    ca_8363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_maxNitr_1727_load_0_ack_1, ack => minSumDecode_CP_6680_elements(340)); -- 
    -- CP-element group 341:  join  transition  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	338 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Sample/rr
      -- 
    rr_8376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(341), ack => ULT_u16_u1_1732_inst_req_0); -- 
    minSumDecode_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(338) & minSumDecode_CP_6680_elements(340);
      gj_minSumDecode_cp_element_group_341 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  transition  input  no-bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_sample_completed_
      -- CP-element group 342: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Sample/ra
      -- 
    ra_8377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u16_u1_1732_inst_ack_0, ack => minSumDecode_CP_6680_elements(342)); -- 
    -- CP-element group 343:  transition  input  no-bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	336 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	26 
    -- CP-element group 343:  members (4) 
      -- CP-element group 343: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/$exit
      -- CP-element group 343: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_update_completed_
      -- CP-element group 343: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_1353/assign_stmt_1725_to_assign_stmt_1733/ULT_u16_u1_1732_Update/ca
      -- 
    ca_8382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ULT_u16_u1_1732_inst_ack_1, ack => minSumDecode_CP_6680_elements(343)); -- 
    -- CP-element group 344:  transition  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	26 
    -- CP-element group 344: successors 
    -- CP-element group 344:  members (1) 
      -- CP-element group 344: 	 branch_block_stmt_1353/if_stmt_1734_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(344) <= minSumDecode_CP_6680_elements(26);
    -- CP-element group 345:  transition  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	26 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_1353/if_stmt_1734_eval_test/$entry
      -- CP-element group 345: 	 branch_block_stmt_1353/if_stmt_1734_eval_test/$exit
      -- CP-element group 345: 	 branch_block_stmt_1353/if_stmt_1734_eval_test/branch_req
      -- 
    branch_req_8390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(345), ack => if_stmt_1734_branch_req_0); -- 
    minSumDecode_CP_6680_elements(345) <= minSumDecode_CP_6680_elements(26);
    -- CP-element group 346:  branch  place  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346: 	349 
    -- CP-element group 346:  members (1) 
      -- CP-element group 346: 	 branch_block_stmt_1353/R_iNsTr_29_1735_place
      -- 
    minSumDecode_CP_6680_elements(346) <= minSumDecode_CP_6680_elements(345);
    -- CP-element group 347:  transition  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (1) 
      -- CP-element group 347: 	 branch_block_stmt_1353/if_stmt_1734_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(347) <= minSumDecode_CP_6680_elements(346);
    -- CP-element group 348:  transition  input  no-bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (2) 
      -- CP-element group 348: 	 branch_block_stmt_1353/if_stmt_1734_if_link/$exit
      -- CP-element group 348: 	 branch_block_stmt_1353/if_stmt_1734_if_link/if_choice_transition
      -- 
    if_choice_transition_8395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1734_branch_ack_1, ack => minSumDecode_CP_6680_elements(348)); -- 
    -- CP-element group 349:  transition  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	346 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (1) 
      -- CP-element group 349: 	 branch_block_stmt_1353/if_stmt_1734_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(349) <= minSumDecode_CP_6680_elements(346);
    -- CP-element group 350:  transition  input  no-bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_1353/if_stmt_1734_else_link/$exit
      -- CP-element group 350: 	 branch_block_stmt_1353/if_stmt_1734_else_link/else_choice_transition
      -- 
    else_choice_transition_8399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1734_branch_ack_0, ack => minSumDecode_CP_6680_elements(350)); -- 
    -- CP-element group 351:  place  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	959 
    -- CP-element group 351:  members (1) 
      -- CP-element group 351: 	 branch_block_stmt_1353/initializeMessagex_xexit_bb_14
      -- 
    minSumDecode_CP_6680_elements(351) <= minSumDecode_CP_6680_elements(348);
    -- CP-element group 352:  place  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	1186 
    -- CP-element group 352:  members (1) 
      -- CP-element group 352: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread
      -- 
    minSumDecode_CP_6680_elements(352) <= minSumDecode_CP_6680_elements(350);
    -- CP-element group 353:  fork  transition  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	27 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (7) 
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/$entry
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_update_start_
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Update/cr
      -- 
    rr_8412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(353), ack => EQ_u16_u1_1745_inst_req_0); -- 
    cr_8417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(353), ack => EQ_u16_u1_1745_inst_req_1); -- 
    minSumDecode_CP_6680_elements(353) <= minSumDecode_CP_6680_elements(27);
    -- CP-element group 354:  transition  input  no-bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Sample/ra
      -- 
    ra_8413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1745_inst_ack_0, ack => minSumDecode_CP_6680_elements(354)); -- 
    -- CP-element group 355:  transition  input  no-bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	28 
    -- CP-element group 355:  members (4) 
      -- CP-element group 355: 	 branch_block_stmt_1353/assign_stmt_1746/$exit
      -- CP-element group 355: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_1353/assign_stmt_1746/EQ_u16_u1_1745_Update/ca
      -- 
    ca_8418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1745_inst_ack_1, ack => minSumDecode_CP_6680_elements(355)); -- 
    -- CP-element group 356:  transition  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	28 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (1) 
      -- CP-element group 356: 	 branch_block_stmt_1353/if_stmt_1747_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(356) <= minSumDecode_CP_6680_elements(28);
    -- CP-element group 357:  transition  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	28 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_1353/if_stmt_1747_eval_test/$entry
      -- CP-element group 357: 	 branch_block_stmt_1353/if_stmt_1747_eval_test/$exit
      -- CP-element group 357: 	 branch_block_stmt_1353/if_stmt_1747_eval_test/branch_req
      -- 
    branch_req_8426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(357), ack => if_stmt_1747_branch_req_0); -- 
    minSumDecode_CP_6680_elements(357) <= minSumDecode_CP_6680_elements(28);
    -- CP-element group 358:  branch  place  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358: 	361 
    -- CP-element group 358:  members (1) 
      -- CP-element group 358: 	 branch_block_stmt_1353/R_iNsTr_40_1748_place
      -- 
    minSumDecode_CP_6680_elements(358) <= minSumDecode_CP_6680_elements(357);
    -- CP-element group 359:  transition  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (1) 
      -- CP-element group 359: 	 branch_block_stmt_1353/if_stmt_1747_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(359) <= minSumDecode_CP_6680_elements(358);
    -- CP-element group 360:  transition  input  no-bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	363 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_1353/if_stmt_1747_if_link/$exit
      -- CP-element group 360: 	 branch_block_stmt_1353/if_stmt_1747_if_link/if_choice_transition
      -- 
    if_choice_transition_8431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1747_branch_ack_1, ack => minSumDecode_CP_6680_elements(360)); -- 
    -- CP-element group 361:  transition  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	358 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (1) 
      -- CP-element group 361: 	 branch_block_stmt_1353/if_stmt_1747_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(361) <= minSumDecode_CP_6680_elements(358);
    -- CP-element group 362:  transition  input  no-bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_1353/if_stmt_1747_else_link/$exit
      -- CP-element group 362: 	 branch_block_stmt_1353/if_stmt_1747_else_link/else_choice_transition
      -- 
    else_choice_transition_8435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1747_branch_ack_0, ack => minSumDecode_CP_6680_elements(362)); -- 
    -- CP-element group 363:  place  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	360 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	978 
    -- CP-element group 363:  members (1) 
      -- CP-element group 363: 	 branch_block_stmt_1353/bb_14_initialize_aPosteriorix_xexit
      -- 
    minSumDecode_CP_6680_elements(363) <= minSumDecode_CP_6680_elements(360);
    -- CP-element group 364:  place  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	962 
    -- CP-element group 364:  members (1) 
      -- CP-element group 364: 	 branch_block_stmt_1353/bb_14_bbx_xnphx_xi18
      -- 
    minSumDecode_CP_6680_elements(364) <= minSumDecode_CP_6680_elements(362);
    -- CP-element group 365:  fork  transition  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	29 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: 	367 
    -- CP-element group 365: 	368 
    -- CP-element group 365: 	369 
    -- CP-element group 365: 	371 
    -- CP-element group 365: 	373 
    -- CP-element group 365: 	376 
    -- CP-element group 365:  members (22) 
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_update_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Update/cr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_update_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Update/cr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_update_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Update/cr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_update_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Update/cr
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_update_start_
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_complete/$entry
      -- CP-element group 365: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_complete/req
      -- 
    rr_8448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => UGT_u16_u1_1758_inst_req_0); -- 
    cr_8453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => UGT_u16_u1_1758_inst_req_1); -- 
    rr_8462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => ADD_u16_u16_1764_inst_req_0); -- 
    cr_8467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => ADD_u16_u16_1764_inst_req_1); -- 
    cr_8481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => type_cast_1768_inst_req_1); -- 
    cr_8495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => ADD_u64_u64_1774_inst_req_1); -- 
    req_8509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(365), ack => MUX_1781_inst_req_1); -- 
    minSumDecode_CP_6680_elements(365) <= minSumDecode_CP_6680_elements(29);
    -- CP-element group 366:  transition  input  no-bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Sample/ra
      -- 
    ra_8449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1758_inst_ack_0, ack => minSumDecode_CP_6680_elements(366)); -- 
    -- CP-element group 367:  transition  input  no-bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	374 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/UGT_u16_u1_1758_Update/ca
      -- 
    ca_8454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1758_inst_ack_1, ack => minSumDecode_CP_6680_elements(367)); -- 
    -- CP-element group 368:  transition  input  no-bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	365 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Sample/ra
      -- 
    ra_8463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1764_inst_ack_0, ack => minSumDecode_CP_6680_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  no-bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u16_u16_1764_Update/ca
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Sample/rr
      -- 
    ca_8468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1764_inst_ack_1, ack => minSumDecode_CP_6680_elements(369)); -- 
    rr_8476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(369), ack => type_cast_1768_inst_req_0); -- 
    -- CP-element group 370:  transition  input  no-bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Sample/ra
      -- 
    ra_8477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_0, ack => minSumDecode_CP_6680_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  no-bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	365 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/type_cast_1768_Update/ca
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Sample/rr
      -- 
    ca_8482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_1, ack => minSumDecode_CP_6680_elements(371)); -- 
    rr_8490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(371), ack => ADD_u64_u64_1774_inst_req_0); -- 
    -- CP-element group 372:  transition  input  no-bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Sample/ra
      -- 
    ra_8491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1774_inst_ack_0, ack => minSumDecode_CP_6680_elements(372)); -- 
    -- CP-element group 373:  transition  input  no-bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	365 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/ADD_u64_u64_1774_Update/ca
      -- 
    ca_8496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1774_inst_ack_1, ack => minSumDecode_CP_6680_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	367 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_start/$entry
      -- CP-element group 374: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_start/req
      -- 
    req_8504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(374), ack => MUX_1781_inst_req_0); -- 
    minSumDecode_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(367) & minSumDecode_CP_6680_elements(373);
      gj_minSumDecode_cp_element_group_374 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  no-bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_start/$exit
      -- CP-element group 375: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_start/ack
      -- 
    ack_8505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1781_inst_ack_0, ack => minSumDecode_CP_6680_elements(375)); -- 
    -- CP-element group 376:  transition  input  no-bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	365 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_complete/$exit
      -- CP-element group 376: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/MUX_1781_complete/ack
      -- 
    ack_8510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1781_inst_ack_1, ack => minSumDecode_CP_6680_elements(376)); -- 
    -- CP-element group 377:  join  transition  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	30 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_1353/assign_stmt_1759_to_assign_stmt_1782/$exit
      -- 
    minSumDecode_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(375) & minSumDecode_CP_6680_elements(376);
      gj_minSumDecode_cp_element_group_377 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	31 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378: 	380 
    -- CP-element group 378: 	381 
    -- CP-element group 378: 	382 
    -- CP-element group 378: 	384 
    -- CP-element group 378: 	387 
    -- CP-element group 378: 	388 
    -- CP-element group 378: 	389 
    -- CP-element group 378: 	391 
    -- CP-element group 378:  members (74) 
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/word_0/cr
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_resize_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_resize_0/index_resize_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_base_plus_offset/sum_rename_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_base_plus_offset/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_complete/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_request/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_base_plus_offset/sum_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_scale_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_resize_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_base_plus_offset/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_scaled_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_complete/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_computed_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_request/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_scale_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_resized_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_scale_0/scale_rename_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_resize_0/index_resize_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_final_index_sum_regn/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/word_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_final_index_sum_regn/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_index_scale_0/scale_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_final_index_sum_regn/ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_final_index_sum_regn/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_root_address_calculated
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_offset_calculated
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_resized_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_scaled_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_computed_0
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_resize_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_resize_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_resize_0/index_resize_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_resize_0/index_resize_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_scale_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_scale_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_scale_0/scale_rename_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_index_scale_0/scale_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_final_index_sum_regn/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_final_index_sum_regn/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_final_index_sum_regn/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_final_index_sum_regn/ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_base_plus_offset/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_base_plus_offset/$exit
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_base_plus_offset/sum_rename_req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1795_base_plus_offset/sum_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_request/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_request/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_complete/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_complete/req
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_root_address_calculated
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/array_obj_ref_1800_offset_calculated
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/word_0/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/word_0/cr
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Update/cr
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Update/cr
      -- 
    req_8551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => addr_of_1796_final_reg_req_1); -- 
    req_8546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => addr_of_1796_final_reg_req_0); -- 
    req_8590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => addr_of_1801_final_reg_req_1); -- 
    req_8585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => addr_of_1801_final_reg_req_0); -- 
    cr_8635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => ptr_deref_1805_load_0_req_1); -- 
    cr_8690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => ptr_deref_1808_store_0_req_1); -- 
    rr_8699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => ADD_u64_u64_1815_inst_req_0); -- 
    cr_8704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => ADD_u64_u64_1815_inst_req_1); -- 
    cr_8718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(378), ack => EQ_u64_u1_1820_inst_req_1); -- 
    minSumDecode_CP_6680_elements(378) <= minSumDecode_CP_6680_elements(31);
    -- CP-element group 379:  transition  input  no-bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	392 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_request/$exit
      -- CP-element group 379: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_request/ack
      -- 
    ack_8547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1796_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(379)); -- 
    -- CP-element group 380:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	383 
    -- CP-element group 380:  members (24) 
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_word_addrgen/$exit
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_word_addrgen/root_register_req
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_word_addrgen/root_register_ack
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/word_0/rr
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_word_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_word_addrgen/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_plus_offset/sum_rename_ack
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_plus_offset/sum_rename_req
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_plus_offset/$exit
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_plus_offset/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_addr_resize/base_resize_ack
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_addr_resize/base_resize_req
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_addr_resize/$exit
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_addr_resize/$entry
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_base_address_resized
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_root_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_complete/$exit
      -- CP-element group 380: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1796_complete/ack
      -- 
    ack_8552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1796_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(380)); -- 
    rr_8624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(380), ack => ptr_deref_1805_load_0_req_0); -- 
    -- CP-element group 381:  transition  input  no-bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	378 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	392 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_request/$exit
      -- CP-element group 381: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_request/ack
      -- CP-element group 381: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_sample_completed_
      -- 
    ack_8586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1801_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(381)); -- 
    -- CP-element group 382:  fork  transition  input  no-bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	378 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	385 
    -- CP-element group 382:  members (19) 
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_complete/$exit
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_word_address_calculated
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_address_calculated
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_address_resized
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_addr_resize/$entry
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_complete/ack
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_addr_resize/$exit
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_addr_resize/base_resize_req
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_root_address_calculated
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/addr_of_1801_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_addr_resize/base_resize_ack
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_plus_offset/$entry
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_plus_offset/$exit
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_plus_offset/sum_rename_req
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_base_plus_offset/sum_rename_ack
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_word_addrgen/$entry
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_word_addrgen/$exit
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_word_addrgen/root_register_req
      -- CP-element group 382: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_word_addrgen/root_register_ack
      -- 
    ack_8591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1801_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(382)); -- 
    -- CP-element group 383:  transition  input  no-bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	380 
    -- CP-element group 383: successors 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/$exit
      -- CP-element group 383: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/word_0/$exit
      -- CP-element group 383: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Sample/word_access_start/word_0/ra
      -- 
    ra_8625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1805_load_0_ack_0, ack => minSumDecode_CP_6680_elements(383)); -- 
    -- CP-element group 384:  transition  input  no-bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	378 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (9) 
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/ptr_deref_1805_Merge/merge_req
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/word_0/ca
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/ptr_deref_1805_Merge/$entry
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/ptr_deref_1805_Merge/$exit
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/ptr_deref_1805_Merge/merge_ack
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/$exit
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1805_Update/word_access_complete/word_0/$exit
      -- 
    ca_8636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1805_load_0_ack_1, ack => minSumDecode_CP_6680_elements(384)); -- 
    -- CP-element group 385:  join  transition  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	382 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (9) 
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/ptr_deref_1808_Split/$entry
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/ptr_deref_1808_Split/$exit
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/ptr_deref_1808_Split/split_req
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/ptr_deref_1808_Split/split_ack
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/$entry
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/word_0/$entry
      -- CP-element group 385: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/word_0/rr
      -- 
    rr_8679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(385), ack => ptr_deref_1808_store_0_req_0); -- 
    minSumDecode_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(382) & minSumDecode_CP_6680_elements(384);
      gj_minSumDecode_cp_element_group_385 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  transition  input  no-bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (5) 
      -- CP-element group 386: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/$exit
      -- CP-element group 386: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/word_0/$exit
      -- CP-element group 386: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Sample/word_access_start/word_0/ra
      -- 
    ra_8680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1808_store_0_ack_0, ack => minSumDecode_CP_6680_elements(386)); -- 
    -- CP-element group 387:  transition  input  no-bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	378 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	392 
    -- CP-element group 387:  members (5) 
      -- CP-element group 387: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/$exit
      -- CP-element group 387: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/word_0/$exit
      -- CP-element group 387: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ptr_deref_1808_Update/word_access_complete/word_0/ca
      -- 
    ca_8691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1808_store_0_ack_1, ack => minSumDecode_CP_6680_elements(387)); -- 
    -- CP-element group 388:  transition  input  no-bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	378 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Sample/ra
      -- 
    ra_8700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1815_inst_ack_0, ack => minSumDecode_CP_6680_elements(388)); -- 
    -- CP-element group 389:  transition  input  output  no-bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	378 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (6) 
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/ADD_u64_u64_1815_Update/ca
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Sample/rr
      -- 
    ca_8705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1815_inst_ack_1, ack => minSumDecode_CP_6680_elements(389)); -- 
    rr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(389), ack => EQ_u64_u1_1820_inst_req_0); -- 
    -- CP-element group 390:  transition  input  no-bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Sample/ra
      -- 
    ra_8714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1820_inst_ack_0, ack => minSumDecode_CP_6680_elements(390)); -- 
    -- CP-element group 391:  transition  input  no-bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	378 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/EQ_u64_u1_1820_Update/ca
      -- 
    ca_8719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1820_inst_ack_1, ack => minSumDecode_CP_6680_elements(391)); -- 
    -- CP-element group 392:  join  transition  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	379 
    -- CP-element group 392: 	381 
    -- CP-element group 392: 	387 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	32 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 branch_block_stmt_1353/assign_stmt_1797_to_assign_stmt_1821/$exit
      -- 
    minSumDecode_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(379) & minSumDecode_CP_6680_elements(381) & minSumDecode_CP_6680_elements(387) & minSumDecode_CP_6680_elements(391);
      gj_minSumDecode_cp_element_group_392 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  transition  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	32 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 branch_block_stmt_1353/if_stmt_1822_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(393) <= minSumDecode_CP_6680_elements(32);
    -- CP-element group 394:  transition  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	32 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_1353/if_stmt_1822_eval_test/$entry
      -- CP-element group 394: 	 branch_block_stmt_1353/if_stmt_1822_eval_test/$exit
      -- CP-element group 394: 	 branch_block_stmt_1353/if_stmt_1822_eval_test/branch_req
      -- 
    branch_req_8727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(394), ack => if_stmt_1822_branch_req_0); -- 
    minSumDecode_CP_6680_elements(394) <= minSumDecode_CP_6680_elements(32);
    -- CP-element group 395:  branch  place  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395: 	398 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 branch_block_stmt_1353/R_exitcond15_1823_place
      -- 
    minSumDecode_CP_6680_elements(395) <= minSumDecode_CP_6680_elements(394);
    -- CP-element group 396:  transition  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 branch_block_stmt_1353/if_stmt_1822_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(396) <= minSumDecode_CP_6680_elements(395);
    -- CP-element group 397:  transition  input  no-bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	400 
    -- CP-element group 397:  members (2) 
      -- CP-element group 397: 	 branch_block_stmt_1353/if_stmt_1822_if_link/$exit
      -- CP-element group 397: 	 branch_block_stmt_1353/if_stmt_1822_if_link/if_choice_transition
      -- 
    if_choice_transition_8732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1822_branch_ack_1, ack => minSumDecode_CP_6680_elements(397)); -- 
    -- CP-element group 398:  transition  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	395 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (1) 
      -- CP-element group 398: 	 branch_block_stmt_1353/if_stmt_1822_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(398) <= minSumDecode_CP_6680_elements(395);
    -- CP-element group 399:  transition  input  no-bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	401 
    -- CP-element group 399:  members (2) 
      -- CP-element group 399: 	 branch_block_stmt_1353/if_stmt_1822_else_link/$exit
      -- CP-element group 399: 	 branch_block_stmt_1353/if_stmt_1822_else_link/else_choice_transition
      -- 
    else_choice_transition_8736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1822_branch_ack_0, ack => minSumDecode_CP_6680_elements(399)); -- 
    -- CP-element group 400:  place  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	397 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	975 
    -- CP-element group 400:  members (1) 
      -- CP-element group 400: 	 branch_block_stmt_1353/bb_16_initialize_aPosteriorix_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(400) <= minSumDecode_CP_6680_elements(397);
    -- CP-element group 401:  place  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	399 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	965 
    -- CP-element group 401:  members (1) 
      -- CP-element group 401: 	 branch_block_stmt_1353/bb_16_bb_16
      -- 
    minSumDecode_CP_6680_elements(401) <= minSumDecode_CP_6680_elements(399);
    -- CP-element group 402:  fork  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	34 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (7) 
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/$entry
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_sample_start_
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_update_start_
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Sample/rr
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Update/cr
      -- 
    rr_8749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(402), ack => EQ_u16_u1_1835_inst_req_0); -- 
    cr_8754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(402), ack => EQ_u16_u1_1835_inst_req_1); -- 
    minSumDecode_CP_6680_elements(402) <= minSumDecode_CP_6680_elements(34);
    -- CP-element group 403:  transition  input  no-bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Sample/ra
      -- 
    ra_8750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1835_inst_ack_0, ack => minSumDecode_CP_6680_elements(403)); -- 
    -- CP-element group 404:  transition  input  no-bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	35 
    -- CP-element group 404:  members (4) 
      -- CP-element group 404: 	 branch_block_stmt_1353/assign_stmt_1836/$exit
      -- CP-element group 404: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_1353/assign_stmt_1836/EQ_u16_u1_1835_Update/ca
      -- 
    ca_8755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1835_inst_ack_1, ack => minSumDecode_CP_6680_elements(404)); -- 
    -- CP-element group 405:  transition  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	35 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (1) 
      -- CP-element group 405: 	 branch_block_stmt_1353/if_stmt_1837_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(405) <= minSumDecode_CP_6680_elements(35);
    -- CP-element group 406:  transition  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	35 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_1353/if_stmt_1837_eval_test/$entry
      -- CP-element group 406: 	 branch_block_stmt_1353/if_stmt_1837_eval_test/$exit
      -- CP-element group 406: 	 branch_block_stmt_1353/if_stmt_1837_eval_test/branch_req
      -- 
    branch_req_8763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(406), ack => if_stmt_1837_branch_req_0); -- 
    minSumDecode_CP_6680_elements(406) <= minSumDecode_CP_6680_elements(35);
    -- CP-element group 407:  branch  place  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407: 	410 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_1353/R_iNsTr_51_1838_place
      -- 
    minSumDecode_CP_6680_elements(407) <= minSumDecode_CP_6680_elements(406);
    -- CP-element group 408:  transition  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (1) 
      -- CP-element group 408: 	 branch_block_stmt_1353/if_stmt_1837_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(408) <= minSumDecode_CP_6680_elements(407);
    -- CP-element group 409:  transition  input  no-bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	412 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_1353/if_stmt_1837_if_link/$exit
      -- CP-element group 409: 	 branch_block_stmt_1353/if_stmt_1837_if_link/if_choice_transition
      -- 
    if_choice_transition_8768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1837_branch_ack_1, ack => minSumDecode_CP_6680_elements(409)); -- 
    -- CP-element group 410:  transition  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	407 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (1) 
      -- CP-element group 410: 	 branch_block_stmt_1353/if_stmt_1837_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(410) <= minSumDecode_CP_6680_elements(407);
    -- CP-element group 411:  transition  input  no-bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	413 
    -- CP-element group 411:  members (2) 
      -- CP-element group 411: 	 branch_block_stmt_1353/if_stmt_1837_else_link/$exit
      -- CP-element group 411: 	 branch_block_stmt_1353/if_stmt_1837_else_link/else_choice_transition
      -- 
    else_choice_transition_8772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1837_branch_ack_0, ack => minSumDecode_CP_6680_elements(411)); -- 
    -- CP-element group 412:  place  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	409 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	999 
    -- CP-element group 412:  members (1) 
      -- CP-element group 412: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_initializeExtrinsicInfox_xexit
      -- 
    minSumDecode_CP_6680_elements(412) <= minSumDecode_CP_6680_elements(409);
    -- CP-element group 413:  place  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	411 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	982 
    -- CP-element group 413:  members (1) 
      -- CP-element group 413: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_bbx_xnphx_xi27
      -- 
    minSumDecode_CP_6680_elements(413) <= minSumDecode_CP_6680_elements(411);
    -- CP-element group 414:  fork  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	36 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414: 	416 
    -- CP-element group 414: 	417 
    -- CP-element group 414: 	418 
    -- CP-element group 414: 	420 
    -- CP-element group 414: 	422 
    -- CP-element group 414: 	425 
    -- CP-element group 414:  members (22) 
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Sample/rr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Sample/rr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Update/cr
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_complete/$entry
      -- CP-element group 414: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_complete/req
      -- 
    rr_8785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => UGT_u16_u1_1848_inst_req_0); -- 
    cr_8790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => UGT_u16_u1_1848_inst_req_1); -- 
    rr_8799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => ADD_u16_u16_1854_inst_req_0); -- 
    cr_8804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => ADD_u16_u16_1854_inst_req_1); -- 
    cr_8818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => type_cast_1858_inst_req_1); -- 
    cr_8832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => ADD_u64_u64_1864_inst_req_1); -- 
    req_8846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(414), ack => MUX_1871_inst_req_1); -- 
    minSumDecode_CP_6680_elements(414) <= minSumDecode_CP_6680_elements(36);
    -- CP-element group 415:  transition  input  no-bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_sample_completed_
      -- CP-element group 415: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Sample/ra
      -- 
    ra_8786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1848_inst_ack_0, ack => minSumDecode_CP_6680_elements(415)); -- 
    -- CP-element group 416:  transition  input  no-bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	423 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/UGT_u16_u1_1848_Update/ca
      -- 
    ca_8791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1848_inst_ack_1, ack => minSumDecode_CP_6680_elements(416)); -- 
    -- CP-element group 417:  transition  input  no-bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	414 
    -- CP-element group 417: successors 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_sample_completed_
      -- CP-element group 417: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Sample/$exit
      -- CP-element group 417: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Sample/ra
      -- 
    ra_8800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1854_inst_ack_0, ack => minSumDecode_CP_6680_elements(417)); -- 
    -- CP-element group 418:  transition  input  output  no-bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	414 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (6) 
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_update_completed_
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Update/$exit
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u16_u16_1854_Update/ca
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Sample/rr
      -- 
    ca_8805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1854_inst_ack_1, ack => minSumDecode_CP_6680_elements(418)); -- 
    rr_8813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(418), ack => type_cast_1858_inst_req_0); -- 
    -- CP-element group 419:  transition  input  no-bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_sample_completed_
      -- CP-element group 419: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Sample/ra
      -- 
    ra_8814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_0, ack => minSumDecode_CP_6680_elements(419)); -- 
    -- CP-element group 420:  transition  input  output  no-bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	414 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (6) 
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/type_cast_1858_Update/ca
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_sample_start_
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Sample/rr
      -- 
    ca_8819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_1, ack => minSumDecode_CP_6680_elements(420)); -- 
    rr_8827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(420), ack => ADD_u64_u64_1864_inst_req_0); -- 
    -- CP-element group 421:  transition  input  no-bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_sample_completed_
      -- CP-element group 421: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Sample/ra
      -- 
    ra_8828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1864_inst_ack_0, ack => minSumDecode_CP_6680_elements(421)); -- 
    -- CP-element group 422:  transition  input  no-bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	414 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_update_completed_
      -- CP-element group 422: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/ADD_u64_u64_1864_Update/ca
      -- 
    ca_8833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1864_inst_ack_1, ack => minSumDecode_CP_6680_elements(422)); -- 
    -- CP-element group 423:  join  transition  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	416 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_sample_start_
      -- CP-element group 423: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_start/$entry
      -- CP-element group 423: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_start/req
      -- 
    req_8841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(423), ack => MUX_1871_inst_req_0); -- 
    minSumDecode_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(416) & minSumDecode_CP_6680_elements(422);
      gj_minSumDecode_cp_element_group_423 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  transition  input  no-bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	426 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_start/$exit
      -- CP-element group 424: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_start/ack
      -- 
    ack_8842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1871_inst_ack_0, ack => minSumDecode_CP_6680_elements(424)); -- 
    -- CP-element group 425:  transition  input  no-bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	414 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_complete/$exit
      -- CP-element group 425: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/MUX_1871_complete/ack
      -- 
    ack_8847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1871_inst_ack_1, ack => minSumDecode_CP_6680_elements(425)); -- 
    -- CP-element group 426:  join  transition  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	424 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	37 
    -- CP-element group 426:  members (1) 
      -- CP-element group 426: 	 branch_block_stmt_1353/assign_stmt_1849_to_assign_stmt_1872/$exit
      -- 
    minSumDecode_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(424) & minSumDecode_CP_6680_elements(425);
      gj_minSumDecode_cp_element_group_426 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  fork  transition  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	38 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427: 	429 
    -- CP-element group 427: 	431 
    -- CP-element group 427: 	432 
    -- CP-element group 427: 	433 
    -- CP-element group 427: 	435 
    -- CP-element group 427:  members (42) 
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_update_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_root_address_calculated
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_offset_calculated
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_resized_0
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_scaled_0
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_computed_0
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_resize_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_resize_0/$exit
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_resize_0/index_resize_req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_resize_0/index_resize_ack
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_scale_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_scale_0/$exit
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_scale_0/scale_rename_req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_index_scale_0/scale_rename_ack
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_final_index_sum_regn/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_final_index_sum_regn/$exit
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_final_index_sum_regn/req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_final_index_sum_regn/ack
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_base_plus_offset/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_base_plus_offset/$exit
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_base_plus_offset/sum_rename_req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/array_obj_ref_1885_base_plus_offset/sum_rename_ack
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_request/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_request/req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_complete/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_complete/req
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_update_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/word_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/word_0/cr
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_update_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Update/cr
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_update_start_
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Update/cr
      -- 
    req_8888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => addr_of_1886_final_reg_req_1); -- 
    req_8883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => addr_of_1886_final_reg_req_0); -- 
    cr_8938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => ptr_deref_1889_store_0_req_1); -- 
    rr_8947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => ADD_u64_u64_1897_inst_req_0); -- 
    cr_8952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => ADD_u64_u64_1897_inst_req_1); -- 
    cr_8966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(427), ack => EQ_u64_u1_1902_inst_req_1); -- 
    minSumDecode_CP_6680_elements(427) <= minSumDecode_CP_6680_elements(38);
    -- CP-element group 428:  transition  input  no-bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	436 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_request/$exit
      -- CP-element group 428: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_request/ack
      -- 
    ack_8884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1886_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(428)); -- 
    -- CP-element group 429:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (28) 
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_complete/$exit
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/addr_of_1886_complete/ack
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_address_calculated
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_word_address_calculated
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_root_address_calculated
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_address_resized
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_addr_resize/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_addr_resize/$exit
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_addr_resize/base_resize_req
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_addr_resize/base_resize_ack
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_plus_offset/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_plus_offset/$exit
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_plus_offset/sum_rename_req
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_base_plus_offset/sum_rename_ack
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_word_addrgen/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_word_addrgen/$exit
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_word_addrgen/root_register_req
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_word_addrgen/root_register_ack
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/ptr_deref_1889_Split/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/ptr_deref_1889_Split/$exit
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/ptr_deref_1889_Split/split_req
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/ptr_deref_1889_Split/split_ack
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/word_0/$entry
      -- CP-element group 429: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/word_0/rr
      -- 
    ack_8889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1886_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(429)); -- 
    rr_8927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(429), ack => ptr_deref_1889_store_0_req_0); -- 
    -- CP-element group 430:  transition  input  no-bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (5) 
      -- CP-element group 430: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_sample_completed_
      -- CP-element group 430: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/$exit
      -- CP-element group 430: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/word_0/$exit
      -- CP-element group 430: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Sample/word_access_start/word_0/ra
      -- 
    ra_8928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1889_store_0_ack_0, ack => minSumDecode_CP_6680_elements(430)); -- 
    -- CP-element group 431:  transition  input  no-bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	427 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	436 
    -- CP-element group 431:  members (5) 
      -- CP-element group 431: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_update_completed_
      -- CP-element group 431: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/$exit
      -- CP-element group 431: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/word_0/$exit
      -- CP-element group 431: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ptr_deref_1889_Update/word_access_complete/word_0/ca
      -- 
    ca_8939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1889_store_0_ack_1, ack => minSumDecode_CP_6680_elements(431)); -- 
    -- CP-element group 432:  transition  input  no-bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	427 
    -- CP-element group 432: successors 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Sample/ra
      -- 
    ra_8948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1897_inst_ack_0, ack => minSumDecode_CP_6680_elements(432)); -- 
    -- CP-element group 433:  transition  input  output  no-bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	427 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (6) 
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/ADD_u64_u64_1897_Update/ca
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Sample/rr
      -- 
    ca_8953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1897_inst_ack_1, ack => minSumDecode_CP_6680_elements(433)); -- 
    rr_8961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(433), ack => EQ_u64_u1_1902_inst_req_0); -- 
    -- CP-element group 434:  transition  input  no-bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_sample_completed_
      -- CP-element group 434: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Sample/ra
      -- 
    ra_8962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1902_inst_ack_0, ack => minSumDecode_CP_6680_elements(434)); -- 
    -- CP-element group 435:  transition  input  no-bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	427 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/EQ_u64_u1_1902_Update/ca
      -- 
    ca_8967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_1902_inst_ack_1, ack => minSumDecode_CP_6680_elements(435)); -- 
    -- CP-element group 436:  join  transition  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	428 
    -- CP-element group 436: 	431 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	39 
    -- CP-element group 436:  members (1) 
      -- CP-element group 436: 	 branch_block_stmt_1353/assign_stmt_1887_to_assign_stmt_1903/$exit
      -- 
    minSumDecode_cp_element_group_436: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_436"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(428) & minSumDecode_CP_6680_elements(431) & minSumDecode_CP_6680_elements(435);
      gj_minSumDecode_cp_element_group_436 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(436), clk => clk, reset => reset); --
    end block;
    -- CP-element group 437:  transition  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	39 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (1) 
      -- CP-element group 437: 	 branch_block_stmt_1353/if_stmt_1904_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(437) <= minSumDecode_CP_6680_elements(39);
    -- CP-element group 438:  transition  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	39 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_1353/if_stmt_1904_eval_test/$entry
      -- CP-element group 438: 	 branch_block_stmt_1353/if_stmt_1904_eval_test/$exit
      -- CP-element group 438: 	 branch_block_stmt_1353/if_stmt_1904_eval_test/branch_req
      -- 
    branch_req_8975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(438), ack => if_stmt_1904_branch_req_0); -- 
    minSumDecode_CP_6680_elements(438) <= minSumDecode_CP_6680_elements(39);
    -- CP-element group 439:  branch  place  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439: 	442 
    -- CP-element group 439:  members (1) 
      -- CP-element group 439: 	 branch_block_stmt_1353/R_exitcond14_1905_place
      -- 
    minSumDecode_CP_6680_elements(439) <= minSumDecode_CP_6680_elements(438);
    -- CP-element group 440:  transition  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (1) 
      -- CP-element group 440: 	 branch_block_stmt_1353/if_stmt_1904_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(440) <= minSumDecode_CP_6680_elements(439);
    -- CP-element group 441:  transition  input  no-bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	444 
    -- CP-element group 441:  members (2) 
      -- CP-element group 441: 	 branch_block_stmt_1353/if_stmt_1904_if_link/$exit
      -- CP-element group 441: 	 branch_block_stmt_1353/if_stmt_1904_if_link/if_choice_transition
      -- 
    if_choice_transition_8980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1904_branch_ack_1, ack => minSumDecode_CP_6680_elements(441)); -- 
    -- CP-element group 442:  transition  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	439 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (1) 
      -- CP-element group 442: 	 branch_block_stmt_1353/if_stmt_1904_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(442) <= minSumDecode_CP_6680_elements(439);
    -- CP-element group 443:  transition  input  no-bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	445 
    -- CP-element group 443:  members (2) 
      -- CP-element group 443: 	 branch_block_stmt_1353/if_stmt_1904_else_link/$exit
      -- CP-element group 443: 	 branch_block_stmt_1353/if_stmt_1904_else_link/else_choice_transition
      -- 
    else_choice_transition_8984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1904_branch_ack_0, ack => minSumDecode_CP_6680_elements(443)); -- 
    -- CP-element group 444:  place  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	441 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	995 
    -- CP-element group 444:  members (1) 
      -- CP-element group 444: 	 branch_block_stmt_1353/bb_20_initializeExtrinsicInfox_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(444) <= minSumDecode_CP_6680_elements(441);
    -- CP-element group 445:  place  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	443 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	985 
    -- CP-element group 445:  members (1) 
      -- CP-element group 445: 	 branch_block_stmt_1353/bb_20_bb_20
      -- 
    minSumDecode_CP_6680_elements(445) <= minSumDecode_CP_6680_elements(443);
    -- CP-element group 446:  fork  transition  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	41 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (7) 
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/$entry
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_sample_start_
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_update_start_
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Sample/crr
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Update/ccr
      -- 
    crr_8997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_8997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(446), ack => call_stmt_1913_call_req_0); -- 
    ccr_9002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_9002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(446), ack => call_stmt_1913_call_req_1); -- 
    minSumDecode_CP_6680_elements(446) <= minSumDecode_CP_6680_elements(41);
    -- CP-element group 447:  transition  input  no-bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Sample/cra
      -- 
    cra_8998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1913_call_ack_0, ack => minSumDecode_CP_6680_elements(447)); -- 
    -- CP-element group 448:  transition  input  no-bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	42 
    -- CP-element group 448:  members (4) 
      -- CP-element group 448: 	 branch_block_stmt_1353/call_stmt_1913/$exit
      -- CP-element group 448: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_1353/call_stmt_1913/call_stmt_1913_Update/cca
      -- 
    cca_9003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1913_call_ack_1, ack => minSumDecode_CP_6680_elements(448)); -- 
    -- CP-element group 449:  fork  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	42 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449: 	451 
    -- CP-element group 449: 	453 
    -- CP-element group 449:  members (16) 
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_update_start_
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_word_address_calculated
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_root_address_calculated
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/word_0/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/word_0/rr
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/word_0/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/word_0/cr
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_update_start_
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Update/cr
      -- 
    cr_9033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(449), ack => LOAD_ncol_ind_1915_load_0_req_1); -- 
    rr_9022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(449), ack => LOAD_ncol_ind_1915_load_0_req_0); -- 
    cr_9052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(449), ack => EQ_u16_u1_1921_inst_req_1); -- 
    minSumDecode_CP_6680_elements(449) <= minSumDecode_CP_6680_elements(42);
    -- CP-element group 450:  transition  input  no-bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450:  members (5) 
      -- CP-element group 450: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/$exit
      -- CP-element group 450: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/word_0/$exit
      -- CP-element group 450: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Sample/word_access_start/word_0/ra
      -- 
    ra_9023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_1915_load_0_ack_0, ack => minSumDecode_CP_6680_elements(450)); -- 
    -- CP-element group 451:  transition  input  output  no-bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (12) 
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_update_completed_
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/$exit
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/word_0/$exit
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/word_access_complete/word_0/ca
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/LOAD_ncol_ind_1915_Merge/$entry
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/LOAD_ncol_ind_1915_Merge/$exit
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/LOAD_ncol_ind_1915_Merge/merge_req
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/LOAD_ncol_ind_1915_Update/LOAD_ncol_ind_1915_Merge/merge_ack
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_sample_start_
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Sample/rr
      -- 
    ca_9034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncol_ind_1915_load_0_ack_1, ack => minSumDecode_CP_6680_elements(451)); -- 
    rr_9047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(451), ack => EQ_u16_u1_1921_inst_req_0); -- 
    -- CP-element group 452:  transition  input  no-bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_sample_completed_
      -- CP-element group 452: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Sample/ra
      -- 
    ra_9048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1921_inst_ack_0, ack => minSumDecode_CP_6680_elements(452)); -- 
    -- CP-element group 453:  transition  input  no-bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	449 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	43 
    -- CP-element group 453:  members (4) 
      -- CP-element group 453: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/$exit
      -- CP-element group 453: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_update_completed_
      -- CP-element group 453: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_1353/assign_stmt_1916_to_assign_stmt_1922/EQ_u16_u1_1921_Update/ca
      -- 
    ca_9053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_1921_inst_ack_1, ack => minSumDecode_CP_6680_elements(453)); -- 
    -- CP-element group 454:  transition  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	43 
    -- CP-element group 454: successors 
    -- CP-element group 454:  members (1) 
      -- CP-element group 454: 	 branch_block_stmt_1353/if_stmt_1923_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(454) <= minSumDecode_CP_6680_elements(43);
    -- CP-element group 455:  transition  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	43 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_1353/if_stmt_1923_eval_test/$entry
      -- CP-element group 455: 	 branch_block_stmt_1353/if_stmt_1923_eval_test/$exit
      -- CP-element group 455: 	 branch_block_stmt_1353/if_stmt_1923_eval_test/branch_req
      -- 
    branch_req_9061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(455), ack => if_stmt_1923_branch_req_0); -- 
    minSumDecode_CP_6680_elements(455) <= minSumDecode_CP_6680_elements(43);
    -- CP-element group 456:  branch  place  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456: 	459 
    -- CP-element group 456:  members (1) 
      -- CP-element group 456: 	 branch_block_stmt_1353/R_iNsTr_67_1924_place
      -- 
    minSumDecode_CP_6680_elements(456) <= minSumDecode_CP_6680_elements(455);
    -- CP-element group 457:  transition  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (1) 
      -- CP-element group 457: 	 branch_block_stmt_1353/if_stmt_1923_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(457) <= minSumDecode_CP_6680_elements(456);
    -- CP-element group 458:  transition  input  no-bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	461 
    -- CP-element group 458:  members (2) 
      -- CP-element group 458: 	 branch_block_stmt_1353/if_stmt_1923_if_link/$exit
      -- CP-element group 458: 	 branch_block_stmt_1353/if_stmt_1923_if_link/if_choice_transition
      -- 
    if_choice_transition_9066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1923_branch_ack_1, ack => minSumDecode_CP_6680_elements(458)); -- 
    -- CP-element group 459:  transition  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	456 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (1) 
      -- CP-element group 459: 	 branch_block_stmt_1353/if_stmt_1923_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(459) <= minSumDecode_CP_6680_elements(456);
    -- CP-element group 460:  transition  input  no-bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	462 
    -- CP-element group 460:  members (2) 
      -- CP-element group 460: 	 branch_block_stmt_1353/if_stmt_1923_else_link/$exit
      -- CP-element group 460: 	 branch_block_stmt_1353/if_stmt_1923_else_link/else_choice_transition
      -- 
    else_choice_transition_9070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1923_branch_ack_0, ack => minSumDecode_CP_6680_elements(460)); -- 
    -- CP-element group 461:  place  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	458 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	1018 
    -- CP-element group 461:  members (1) 
      -- CP-element group 461: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_update_aPosteriorix_xexit
      -- 
    minSumDecode_CP_6680_elements(461) <= minSumDecode_CP_6680_elements(458);
    -- CP-element group 462:  place  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	460 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	1002 
    -- CP-element group 462:  members (1) 
      -- CP-element group 462: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_bbx_xnphx_xi54
      -- 
    minSumDecode_CP_6680_elements(462) <= minSumDecode_CP_6680_elements(460);
    -- CP-element group 463:  fork  transition  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	44 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463: 	465 
    -- CP-element group 463: 	466 
    -- CP-element group 463: 	467 
    -- CP-element group 463: 	469 
    -- CP-element group 463: 	471 
    -- CP-element group 463: 	474 
    -- CP-element group 463:  members (22) 
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_update_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Sample/rr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Update/cr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_update_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Sample/rr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Update/cr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_update_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Update/cr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_update_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Update/cr
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_update_start_
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_complete/$entry
      -- CP-element group 463: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_complete/req
      -- 
    rr_9083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => UGT_u16_u1_1934_inst_req_0); -- 
    cr_9088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => UGT_u16_u1_1934_inst_req_1); -- 
    rr_9097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => ADD_u16_u16_1940_inst_req_0); -- 
    cr_9102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => ADD_u16_u16_1940_inst_req_1); -- 
    cr_9116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => type_cast_1944_inst_req_1); -- 
    cr_9130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => ADD_u64_u64_1950_inst_req_1); -- 
    req_9144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(463), ack => MUX_1957_inst_req_1); -- 
    minSumDecode_CP_6680_elements(463) <= minSumDecode_CP_6680_elements(44);
    -- CP-element group 464:  transition  input  no-bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Sample/ra
      -- 
    ra_9084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1934_inst_ack_0, ack => minSumDecode_CP_6680_elements(464)); -- 
    -- CP-element group 465:  transition  input  no-bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	463 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	472 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/UGT_u16_u1_1934_Update/ca
      -- 
    ca_9089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_1934_inst_ack_1, ack => minSumDecode_CP_6680_elements(465)); -- 
    -- CP-element group 466:  transition  input  no-bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	463 
    -- CP-element group 466: successors 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_sample_completed_
      -- CP-element group 466: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Sample/$exit
      -- CP-element group 466: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Sample/ra
      -- 
    ra_9098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1940_inst_ack_0, ack => minSumDecode_CP_6680_elements(466)); -- 
    -- CP-element group 467:  transition  input  output  no-bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	463 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467:  members (6) 
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_update_completed_
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Update/$exit
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u16_u16_1940_Update/ca
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_sample_start_
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Sample/$entry
      -- CP-element group 467: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Sample/rr
      -- 
    ca_9103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1940_inst_ack_1, ack => minSumDecode_CP_6680_elements(467)); -- 
    rr_9111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(467), ack => type_cast_1944_inst_req_0); -- 
    -- CP-element group 468:  transition  input  no-bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Sample/ra
      -- 
    ra_9112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_0, ack => minSumDecode_CP_6680_elements(468)); -- 
    -- CP-element group 469:  transition  input  output  no-bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	463 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	470 
    -- CP-element group 469:  members (6) 
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/type_cast_1944_Update/ca
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Sample/rr
      -- 
    ca_9117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_1, ack => minSumDecode_CP_6680_elements(469)); -- 
    rr_9125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(469), ack => ADD_u64_u64_1950_inst_req_0); -- 
    -- CP-element group 470:  transition  input  no-bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	469 
    -- CP-element group 470: successors 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_sample_completed_
      -- CP-element group 470: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Sample/$exit
      -- CP-element group 470: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Sample/ra
      -- 
    ra_9126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1950_inst_ack_0, ack => minSumDecode_CP_6680_elements(470)); -- 
    -- CP-element group 471:  transition  input  no-bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	463 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_update_completed_
      -- CP-element group 471: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Update/$exit
      -- CP-element group 471: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/ADD_u64_u64_1950_Update/ca
      -- 
    ca_9131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1950_inst_ack_1, ack => minSumDecode_CP_6680_elements(471)); -- 
    -- CP-element group 472:  join  transition  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	465 
    -- CP-element group 472: 	471 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_sample_start_
      -- CP-element group 472: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_start/$entry
      -- CP-element group 472: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_start/req
      -- 
    req_9139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(472), ack => MUX_1957_inst_req_0); -- 
    minSumDecode_cp_element_group_472: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_472"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(465) & minSumDecode_CP_6680_elements(471);
      gj_minSumDecode_cp_element_group_472 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(472), clk => clk, reset => reset); --
    end block;
    -- CP-element group 473:  transition  input  no-bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	475 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_sample_completed_
      -- CP-element group 473: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_start/$exit
      -- CP-element group 473: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_start/ack
      -- 
    ack_9140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1957_inst_ack_0, ack => minSumDecode_CP_6680_elements(473)); -- 
    -- CP-element group 474:  transition  input  no-bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	463 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_update_completed_
      -- CP-element group 474: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_complete/$exit
      -- CP-element group 474: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/MUX_1957_complete/ack
      -- 
    ack_9145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1957_inst_ack_1, ack => minSumDecode_CP_6680_elements(474)); -- 
    -- CP-element group 475:  join  transition  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	473 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	45 
    -- CP-element group 475:  members (1) 
      -- CP-element group 475: 	 branch_block_stmt_1353/assign_stmt_1935_to_assign_stmt_1958/$exit
      -- 
    minSumDecode_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(473) & minSumDecode_CP_6680_elements(474);
      gj_minSumDecode_cp_element_group_475 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  fork  transition  output  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	46 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	477 
    -- CP-element group 476: 	478 
    -- CP-element group 476: 	479 
    -- CP-element group 476: 	480 
    -- CP-element group 476: 	482 
    -- CP-element group 476: 	484 
    -- CP-element group 476: 	486 
    -- CP-element group 476: 	488 
    -- CP-element group 476: 	490 
    -- CP-element group 476: 	492 
    -- CP-element group 476: 	494 
    -- CP-element group 476: 	497 
    -- CP-element group 476: 	500 
    -- CP-element group 476: 	501 
    -- CP-element group 476: 	502 
    -- CP-element group 476: 	504 
    -- CP-element group 476:  members (78) 
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_sample_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_root_address_calculated
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_offset_calculated
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_resized_0
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_scaled_0
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_computed_0
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_resize_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_resize_0/$exit
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_resize_0/index_resize_req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_resize_0/index_resize_ack
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_scale_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_scale_0/$exit
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_scale_0/scale_rename_req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_index_scale_0/scale_rename_ack
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_final_index_sum_regn/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_final_index_sum_regn/$exit
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_final_index_sum_regn/req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_final_index_sum_regn/ack
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_base_plus_offset/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_base_plus_offset/$exit
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_base_plus_offset/sum_rename_req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1971_base_plus_offset/sum_rename_ack
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_request/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_request/req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_complete/req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_sample_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Sample/rr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_complete/req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_complete/req
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_sample_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_update_start_
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Sample/rr
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Update/cr
      -- 
    req_9186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => addr_of_1972_final_reg_req_1); -- 
    req_9181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => addr_of_1972_final_reg_req_0); -- 
    rr_9195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_u64_u64_1978_inst_req_0); -- 
    cr_9200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_u64_u64_1978_inst_req_1); -- 
    req_9239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => addr_of_1983_final_reg_req_1); -- 
    cr_9284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ptr_deref_1987_load_0_req_1); -- 
    cr_9303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_u16_u16_1993_inst_req_1); -- 
    cr_9348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ptr_deref_1997_load_0_req_1); -- 
    cr_9367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => type_cast_2001_inst_req_1); -- 
    req_9406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => addr_of_2006_final_reg_req_1); -- 
    cr_9451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ptr_deref_2010_load_0_req_1); -- 
    cr_9470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_f32_f32_2015_inst_req_1); -- 
    cr_9520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ptr_deref_2018_store_0_req_1); -- 
    rr_9529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_u64_u64_2025_inst_req_0); -- 
    cr_9534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => ADD_u64_u64_2025_inst_req_1); -- 
    cr_9548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(476), ack => EQ_u64_u1_2030_inst_req_1); -- 
    minSumDecode_CP_6680_elements(476) <= minSumDecode_CP_6680_elements(46);
    -- CP-element group 477:  transition  input  no-bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	476 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	506 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_sample_completed_
      -- CP-element group 477: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_request/$exit
      -- CP-element group 477: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_request/ack
      -- 
    ack_9182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1972_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(477)); -- 
    -- CP-element group 478:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	476 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	487 
    -- CP-element group 478:  members (24) 
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_update_completed_
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_complete/$exit
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1972_complete/ack
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_sample_start_
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_address_calculated
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_word_address_calculated
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_root_address_calculated
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_address_resized
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_addr_resize/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_addr_resize/$exit
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_addr_resize/base_resize_req
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_addr_resize/base_resize_ack
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_plus_offset/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_plus_offset/$exit
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_plus_offset/sum_rename_req
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_base_plus_offset/sum_rename_ack
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_word_addrgen/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_word_addrgen/$exit
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_word_addrgen/root_register_req
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_word_addrgen/root_register_ack
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/word_0/$entry
      -- CP-element group 478: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/word_0/rr
      -- 
    ack_9187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1972_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(478)); -- 
    rr_9337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(478), ack => ptr_deref_1997_load_0_req_0); -- 
    -- CP-element group 479:  transition  input  no-bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	476 
    -- CP-element group 479: successors 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_sample_completed_
      -- CP-element group 479: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Sample/$exit
      -- CP-element group 479: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Sample/ra
      -- 
    ra_9196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1978_inst_ack_0, ack => minSumDecode_CP_6680_elements(479)); -- 
    -- CP-element group 480:  transition  input  output  no-bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	476 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (27) 
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_update_completed_
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Update/$exit
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_1978_Update/ca
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_sample_start_
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_root_address_calculated
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_offset_calculated
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_resized_0
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_scaled_0
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_computed_0
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_resize_0/$entry
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_resize_0/$exit
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_resize_0/index_resize_req
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_resize_0/index_resize_ack
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_scale_0/$entry
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_scale_0/$exit
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_scale_0/scale_rename_req
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_index_scale_0/scale_rename_ack
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_final_index_sum_regn/$entry
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_final_index_sum_regn/$exit
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_final_index_sum_regn/req
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_final_index_sum_regn/ack
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_base_plus_offset/$entry
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_base_plus_offset/$exit
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_base_plus_offset/sum_rename_req
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_1982_base_plus_offset/sum_rename_ack
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_request/$entry
      -- CP-element group 480: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_request/req
      -- 
    ca_9201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1978_inst_ack_1, ack => minSumDecode_CP_6680_elements(480)); -- 
    req_9234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(480), ack => addr_of_1983_final_reg_req_0); -- 
    -- CP-element group 481:  transition  input  no-bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	506 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_sample_completed_
      -- CP-element group 481: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_request/$exit
      -- CP-element group 481: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_request/ack
      -- 
    ack_9235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(481)); -- 
    -- CP-element group 482:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	476 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482:  members (24) 
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_complete/$exit
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_1983_complete/ack
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_word_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_root_address_calculated
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_address_resized
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_addr_resize/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_addr_resize/$exit
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_addr_resize/base_resize_req
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_addr_resize/base_resize_ack
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_plus_offset/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_plus_offset/$exit
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_plus_offset/sum_rename_req
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_base_plus_offset/sum_rename_ack
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_word_addrgen/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_word_addrgen/$exit
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_word_addrgen/root_register_req
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_word_addrgen/root_register_ack
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/word_0/rr
      -- 
    ack_9240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1983_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(482)); -- 
    rr_9273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(482), ack => ptr_deref_1987_load_0_req_0); -- 
    -- CP-element group 483:  transition  input  no-bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483:  members (5) 
      -- CP-element group 483: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_sample_completed_
      -- CP-element group 483: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/$exit
      -- CP-element group 483: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/word_0/$exit
      -- CP-element group 483: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Sample/word_access_start/word_0/ra
      -- 
    ra_9274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1987_load_0_ack_0, ack => minSumDecode_CP_6680_elements(483)); -- 
    -- CP-element group 484:  transition  input  output  no-bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	476 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (12) 
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_update_completed_
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/$exit
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/word_0/$exit
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/word_access_complete/word_0/ca
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/ptr_deref_1987_Merge/$entry
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/ptr_deref_1987_Merge/$exit
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/ptr_deref_1987_Merge/merge_req
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1987_Update/ptr_deref_1987_Merge/merge_ack
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_sample_start_
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Sample/rr
      -- 
    ca_9285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1987_load_0_ack_1, ack => minSumDecode_CP_6680_elements(484)); -- 
    rr_9298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(484), ack => ADD_u16_u16_1993_inst_req_0); -- 
    -- CP-element group 485:  transition  input  no-bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_sample_completed_
      -- CP-element group 485: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Sample/ra
      -- 
    ra_9299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1993_inst_ack_0, ack => minSumDecode_CP_6680_elements(485)); -- 
    -- CP-element group 486:  transition  input  output  no-bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	476 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	489 
    -- CP-element group 486:  members (6) 
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_update_completed_
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u16_u16_1993_Update/ca
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Sample/rr
      -- 
    ca_9304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1993_inst_ack_1, ack => minSumDecode_CP_6680_elements(486)); -- 
    rr_9362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(486), ack => type_cast_2001_inst_req_0); -- 
    -- CP-element group 487:  transition  input  no-bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	478 
    -- CP-element group 487: successors 
    -- CP-element group 487:  members (5) 
      -- CP-element group 487: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/$exit
      -- CP-element group 487: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/word_0/$exit
      -- CP-element group 487: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Sample/word_access_start/word_0/ra
      -- 
    ra_9338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1997_load_0_ack_0, ack => minSumDecode_CP_6680_elements(487)); -- 
    -- CP-element group 488:  transition  input  no-bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	476 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	495 
    -- CP-element group 488:  members (9) 
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/$exit
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/word_0/$exit
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/word_access_complete/word_0/ca
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/ptr_deref_1997_Merge/$entry
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/ptr_deref_1997_Merge/$exit
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/ptr_deref_1997_Merge/merge_req
      -- CP-element group 488: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_1997_Update/ptr_deref_1997_Merge/merge_ack
      -- 
    ca_9349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1997_load_0_ack_1, ack => minSumDecode_CP_6680_elements(488)); -- 
    -- CP-element group 489:  transition  input  no-bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	486 
    -- CP-element group 489: successors 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Sample/ra
      -- 
    ra_9363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_0, ack => minSumDecode_CP_6680_elements(489)); -- 
    -- CP-element group 490:  transition  input  output  no-bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	476 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (27) 
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/type_cast_2001_Update/ca
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_root_address_calculated
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_offset_calculated
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_resized_0
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_scaled_0
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_computed_0
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_resize_0/$entry
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_resize_0/$exit
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_resize_0/index_resize_req
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_resize_0/index_resize_ack
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_scale_0/$entry
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_scale_0/$exit
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_scale_0/scale_rename_req
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_index_scale_0/scale_rename_ack
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_final_index_sum_regn/$entry
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_final_index_sum_regn/$exit
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_final_index_sum_regn/req
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_final_index_sum_regn/ack
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_base_plus_offset/$entry
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_base_plus_offset/$exit
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_base_plus_offset/sum_rename_req
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/array_obj_ref_2005_base_plus_offset/sum_rename_ack
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_request/$entry
      -- CP-element group 490: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_request/req
      -- 
    ca_9368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2001_inst_ack_1, ack => minSumDecode_CP_6680_elements(490)); -- 
    req_9401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(490), ack => addr_of_2006_final_reg_req_0); -- 
    -- CP-element group 491:  transition  input  no-bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	506 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_request/$exit
      -- CP-element group 491: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_request/ack
      -- 
    ack_9402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2006_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(491)); -- 
    -- CP-element group 492:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	476 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492: 	498 
    -- CP-element group 492:  members (40) 
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_complete/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/addr_of_2006_complete/ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_sample_start_
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_word_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_root_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_address_resized
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_addr_resize/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_addr_resize/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_addr_resize/base_resize_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_addr_resize/base_resize_ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_plus_offset/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_plus_offset/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_plus_offset/sum_rename_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_base_plus_offset/sum_rename_ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_word_addrgen/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_word_addrgen/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_word_addrgen/root_register_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_word_addrgen/root_register_ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/word_0/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/word_0/rr
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_word_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_root_address_calculated
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_address_resized
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_addr_resize/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_addr_resize/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_addr_resize/base_resize_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_addr_resize/base_resize_ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_plus_offset/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_plus_offset/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_plus_offset/sum_rename_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_base_plus_offset/sum_rename_ack
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_word_addrgen/$entry
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_word_addrgen/$exit
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_word_addrgen/root_register_req
      -- CP-element group 492: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_word_addrgen/root_register_ack
      -- 
    ack_9407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2006_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(492)); -- 
    rr_9440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(492), ack => ptr_deref_2010_load_0_req_0); -- 
    -- CP-element group 493:  transition  input  no-bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	505 
    -- CP-element group 493:  members (5) 
      -- CP-element group 493: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_sample_completed_
      -- CP-element group 493: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/$exit
      -- CP-element group 493: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/$exit
      -- CP-element group 493: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/word_0/$exit
      -- CP-element group 493: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Sample/word_access_start/word_0/ra
      -- 
    ra_9441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2010_load_0_ack_0, ack => minSumDecode_CP_6680_elements(493)); -- 
    -- CP-element group 494:  transition  input  no-bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	476 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (9) 
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_update_completed_
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/$exit
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/$exit
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/word_0/$exit
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/word_access_complete/word_0/ca
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/ptr_deref_2010_Merge/$entry
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/ptr_deref_2010_Merge/$exit
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/ptr_deref_2010_Merge/merge_req
      -- CP-element group 494: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_Update/ptr_deref_2010_Merge/merge_ack
      -- 
    ca_9452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2010_load_0_ack_1, ack => minSumDecode_CP_6680_elements(494)); -- 
    -- CP-element group 495:  join  transition  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	488 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_sample_start_
      -- CP-element group 495: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Sample/rr
      -- 
    rr_9465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(495), ack => ADD_f32_f32_2015_inst_req_0); -- 
    minSumDecode_cp_element_group_495: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_495"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(488) & minSumDecode_CP_6680_elements(494);
      gj_minSumDecode_cp_element_group_495 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(495), clk => clk, reset => reset); --
    end block;
    -- CP-element group 496:  transition  input  no-bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_sample_completed_
      -- CP-element group 496: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Sample/$exit
      -- CP-element group 496: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Sample/ra
      -- 
    ra_9466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2015_inst_ack_0, ack => minSumDecode_CP_6680_elements(496)); -- 
    -- CP-element group 497:  transition  input  no-bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	476 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_update_completed_
      -- CP-element group 497: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Update/$exit
      -- CP-element group 497: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_f32_f32_2015_Update/ca
      -- 
    ca_9471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_f32_f32_2015_inst_ack_1, ack => minSumDecode_CP_6680_elements(497)); -- 
    -- CP-element group 498:  join  transition  output  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	492 
    -- CP-element group 498: 	497 
    -- CP-element group 498: 	505 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498:  members (9) 
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_sample_start_
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/ptr_deref_2018_Split/$entry
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/ptr_deref_2018_Split/$exit
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/ptr_deref_2018_Split/split_req
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/ptr_deref_2018_Split/split_ack
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/$entry
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/word_0/$entry
      -- CP-element group 498: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/word_0/rr
      -- 
    rr_9509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(498), ack => ptr_deref_2018_store_0_req_0); -- 
    minSumDecode_cp_element_group_498: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_498"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(492) & minSumDecode_CP_6680_elements(497) & minSumDecode_CP_6680_elements(505);
      gj_minSumDecode_cp_element_group_498 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 499:  transition  input  no-bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	498 
    -- CP-element group 499: successors 
    -- CP-element group 499:  members (5) 
      -- CP-element group 499: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_sample_completed_
      -- CP-element group 499: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/$exit
      -- CP-element group 499: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/$exit
      -- CP-element group 499: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/word_0/$exit
      -- CP-element group 499: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Sample/word_access_start/word_0/ra
      -- 
    ra_9510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_0_ack_0, ack => minSumDecode_CP_6680_elements(499)); -- 
    -- CP-element group 500:  transition  input  no-bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	476 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	506 
    -- CP-element group 500:  members (5) 
      -- CP-element group 500: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_update_completed_
      -- CP-element group 500: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/$exit
      -- CP-element group 500: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/$exit
      -- CP-element group 500: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/word_0/$exit
      -- CP-element group 500: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2018_Update/word_access_complete/word_0/ca
      -- 
    ca_9521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2018_store_0_ack_1, ack => minSumDecode_CP_6680_elements(500)); -- 
    -- CP-element group 501:  transition  input  no-bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	476 
    -- CP-element group 501: successors 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Sample/ra
      -- 
    ra_9530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2025_inst_ack_0, ack => minSumDecode_CP_6680_elements(501)); -- 
    -- CP-element group 502:  transition  input  output  no-bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	476 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502:  members (6) 
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Sample/$entry
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Sample/rr
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ADD_u64_u64_2025_Update/ca
      -- CP-element group 502: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_sample_start_
      -- 
    ca_9535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2025_inst_ack_1, ack => minSumDecode_CP_6680_elements(502)); -- 
    rr_9543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(502), ack => EQ_u64_u1_2030_inst_req_0); -- 
    -- CP-element group 503:  transition  input  no-bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: successors 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Sample/ra
      -- CP-element group 503: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Sample/$exit
      -- CP-element group 503: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_sample_completed_
      -- 
    ra_9544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2030_inst_ack_0, ack => minSumDecode_CP_6680_elements(503)); -- 
    -- CP-element group 504:  transition  input  no-bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	476 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	506 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Update/ca
      -- CP-element group 504: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_Update/$exit
      -- CP-element group 504: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/EQ_u64_u1_2030_update_completed_
      -- 
    ca_9549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2030_inst_ack_1, ack => minSumDecode_CP_6680_elements(504)); -- 
    -- CP-element group 505:  transition  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	493 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	498 
    -- CP-element group 505:  members (1) 
      -- CP-element group 505: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/ptr_deref_2010_ptr_deref_2018_delay
      -- 
    -- Element group minSumDecode_CP_6680_elements(505) is a control-delay.
    cp_element_505_delay: control_delay_element  generic map(name => " 505_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(493), ack => minSumDecode_CP_6680_elements(505), clk => clk, reset =>reset);
    -- CP-element group 506:  join  transition  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	477 
    -- CP-element group 506: 	481 
    -- CP-element group 506: 	491 
    -- CP-element group 506: 	500 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	47 
    -- CP-element group 506:  members (1) 
      -- CP-element group 506: 	 branch_block_stmt_1353/assign_stmt_1973_to_assign_stmt_2031/$exit
      -- 
    minSumDecode_cp_element_group_506: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_506"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(477) & minSumDecode_CP_6680_elements(481) & minSumDecode_CP_6680_elements(491) & minSumDecode_CP_6680_elements(500) & minSumDecode_CP_6680_elements(504);
      gj_minSumDecode_cp_element_group_506 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(506), clk => clk, reset => reset); --
    end block;
    -- CP-element group 507:  transition  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	47 
    -- CP-element group 507: successors 
    -- CP-element group 507:  members (1) 
      -- CP-element group 507: 	 branch_block_stmt_1353/if_stmt_2032_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(507) <= minSumDecode_CP_6680_elements(47);
    -- CP-element group 508:  transition  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	47 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	509 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_1353/if_stmt_2032_eval_test/$exit
      -- CP-element group 508: 	 branch_block_stmt_1353/if_stmt_2032_eval_test/$entry
      -- CP-element group 508: 	 branch_block_stmt_1353/if_stmt_2032_eval_test/branch_req
      -- 
    branch_req_9558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(508), ack => if_stmt_2032_branch_req_0); -- 
    minSumDecode_CP_6680_elements(508) <= minSumDecode_CP_6680_elements(47);
    -- CP-element group 509:  branch  place  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	508 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	510 
    -- CP-element group 509: 	512 
    -- CP-element group 509:  members (1) 
      -- CP-element group 509: 	 branch_block_stmt_1353/R_exitcond12_2033_place
      -- 
    minSumDecode_CP_6680_elements(509) <= minSumDecode_CP_6680_elements(508);
    -- CP-element group 510:  transition  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	509 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	511 
    -- CP-element group 510:  members (1) 
      -- CP-element group 510: 	 branch_block_stmt_1353/if_stmt_2032_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(510) <= minSumDecode_CP_6680_elements(509);
    -- CP-element group 511:  transition  input  no-bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	510 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	514 
    -- CP-element group 511:  members (2) 
      -- CP-element group 511: 	 branch_block_stmt_1353/if_stmt_2032_if_link/if_choice_transition
      -- CP-element group 511: 	 branch_block_stmt_1353/if_stmt_2032_if_link/$exit
      -- 
    if_choice_transition_9563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2032_branch_ack_1, ack => minSumDecode_CP_6680_elements(511)); -- 
    -- CP-element group 512:  transition  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	509 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	513 
    -- CP-element group 512:  members (1) 
      -- CP-element group 512: 	 branch_block_stmt_1353/if_stmt_2032_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(512) <= minSumDecode_CP_6680_elements(509);
    -- CP-element group 513:  transition  input  no-bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	512 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	515 
    -- CP-element group 513:  members (2) 
      -- CP-element group 513: 	 branch_block_stmt_1353/if_stmt_2032_else_link/else_choice_transition
      -- CP-element group 513: 	 branch_block_stmt_1353/if_stmt_2032_else_link/$exit
      -- 
    else_choice_transition_9567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2032_branch_ack_0, ack => minSumDecode_CP_6680_elements(513)); -- 
    -- CP-element group 514:  place  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	511 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	1015 
    -- CP-element group 514:  members (1) 
      -- CP-element group 514: 	 branch_block_stmt_1353/bb_24_update_aPosteriorix_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(514) <= minSumDecode_CP_6680_elements(511);
    -- CP-element group 515:  place  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	513 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	1005 
    -- CP-element group 515:  members (1) 
      -- CP-element group 515: 	 branch_block_stmt_1353/bb_24_bb_24
      -- 
    minSumDecode_CP_6680_elements(515) <= minSumDecode_CP_6680_elements(513);
    -- CP-element group 516:  fork  transition  output  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	49 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	517 
    -- CP-element group 516: 	518 
    -- CP-element group 516: 	519 
    -- CP-element group 516: 	520 
    -- CP-element group 516: 	522 
    -- CP-element group 516:  members (32) 
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_update_start_
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_word_address_calculated
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_root_address_calculated
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/word_0/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/word_0/rr
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/word_0/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_sample_start_
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/word_0/cr
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/word_0/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/word_0/rr
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/word_0/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Update/cr
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/STORE_is_decoded_2041_Split/split_ack
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/STORE_is_decoded_2041_Split/split_req
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/STORE_is_decoded_2041_Split/$exit
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/STORE_is_decoded_2041_Split/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_root_address_calculated
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_word_address_calculated
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_update_start_
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_update_start_
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_sample_start_
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/$entry
      -- CP-element group 516: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/word_0/cr
      -- 
    cr_9604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(516), ack => STORE_is_decoded_2041_store_0_req_1); -- 
    rr_9593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(516), ack => STORE_is_decoded_2041_store_0_req_0); -- 
    cr_9632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(516), ack => LOAD_ncols_2046_load_0_req_1); -- 
    rr_9621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(516), ack => LOAD_ncols_2046_load_0_req_0); -- 
    cr_9651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(516), ack => EQ_u16_u1_2052_inst_req_1); -- 
    minSumDecode_CP_6680_elements(516) <= minSumDecode_CP_6680_elements(49);
    -- CP-element group 517:  transition  input  no-bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	516 
    -- CP-element group 517: successors 
    -- CP-element group 517:  members (5) 
      -- CP-element group 517: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/word_0/ra
      -- CP-element group 517: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/word_0/$exit
      -- CP-element group 517: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/word_access_start/$exit
      -- CP-element group 517: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_sample_completed_
      -- 
    ra_9594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2041_store_0_ack_0, ack => minSumDecode_CP_6680_elements(517)); -- 
    -- CP-element group 518:  transition  input  no-bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	516 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	523 
    -- CP-element group 518:  members (5) 
      -- CP-element group 518: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/word_0/ca
      -- CP-element group 518: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/word_0/$exit
      -- CP-element group 518: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/word_access_complete/$exit
      -- CP-element group 518: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_Update/$exit
      -- CP-element group 518: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/STORE_is_decoded_2041_update_completed_
      -- 
    ca_9605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2041_store_0_ack_1, ack => minSumDecode_CP_6680_elements(518)); -- 
    -- CP-element group 519:  transition  input  no-bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	516 
    -- CP-element group 519: successors 
    -- CP-element group 519:  members (5) 
      -- CP-element group 519: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/$exit
      -- CP-element group 519: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/$exit
      -- CP-element group 519: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/word_0/$exit
      -- CP-element group 519: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Sample/word_access_start/word_0/ra
      -- CP-element group 519: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_sample_completed_
      -- 
    ra_9622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_2046_load_0_ack_0, ack => minSumDecode_CP_6680_elements(519)); -- 
    -- CP-element group 520:  transition  input  output  no-bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	516 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	521 
    -- CP-element group 520:  members (12) 
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_update_completed_
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/$exit
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/$exit
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Sample/rr
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Sample/$entry
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_sample_start_
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/LOAD_ncols_2046_Merge/merge_ack
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/LOAD_ncols_2046_Merge/merge_req
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/LOAD_ncols_2046_Merge/$exit
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/LOAD_ncols_2046_Merge/$entry
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/word_0/ca
      -- CP-element group 520: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/LOAD_ncols_2046_Update/word_access_complete/word_0/$exit
      -- 
    ca_9633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_2046_load_0_ack_1, ack => minSumDecode_CP_6680_elements(520)); -- 
    rr_9646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(520), ack => EQ_u16_u1_2052_inst_req_0); -- 
    -- CP-element group 521:  transition  input  no-bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	520 
    -- CP-element group 521: successors 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_sample_completed_
      -- CP-element group 521: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Sample/ra
      -- CP-element group 521: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Sample/$exit
      -- 
    ra_9647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2052_inst_ack_0, ack => minSumDecode_CP_6680_elements(521)); -- 
    -- CP-element group 522:  transition  input  no-bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	516 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	523 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Update/ca
      -- CP-element group 522: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_Update/$exit
      -- CP-element group 522: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/EQ_u16_u1_2052_update_completed_
      -- 
    ca_9652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2052_inst_ack_1, ack => minSumDecode_CP_6680_elements(522)); -- 
    -- CP-element group 523:  join  transition  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	518 
    -- CP-element group 523: 	522 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	50 
    -- CP-element group 523:  members (1) 
      -- CP-element group 523: 	 branch_block_stmt_1353/assign_stmt_2044_to_assign_stmt_2053/$exit
      -- 
    minSumDecode_cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(518) & minSumDecode_CP_6680_elements(522);
      gj_minSumDecode_cp_element_group_523 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 524:  transition  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	50 
    -- CP-element group 524: successors 
    -- CP-element group 524:  members (1) 
      -- CP-element group 524: 	 branch_block_stmt_1353/if_stmt_2054_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(524) <= minSumDecode_CP_6680_elements(50);
    -- CP-element group 525:  transition  output  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	50 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_1353/if_stmt_2054_eval_test/branch_req
      -- CP-element group 525: 	 branch_block_stmt_1353/if_stmt_2054_eval_test/$exit
      -- CP-element group 525: 	 branch_block_stmt_1353/if_stmt_2054_eval_test/$entry
      -- 
    branch_req_9660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(525), ack => if_stmt_2054_branch_req_0); -- 
    minSumDecode_CP_6680_elements(525) <= minSumDecode_CP_6680_elements(50);
    -- CP-element group 526:  branch  place  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	525 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526: 	529 
    -- CP-element group 526:  members (1) 
      -- CP-element group 526: 	 branch_block_stmt_1353/R_iNsTr_84_2055_place
      -- 
    minSumDecode_CP_6680_elements(526) <= minSumDecode_CP_6680_elements(525);
    -- CP-element group 527:  transition  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	528 
    -- CP-element group 527:  members (1) 
      -- CP-element group 527: 	 branch_block_stmt_1353/if_stmt_2054_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(527) <= minSumDecode_CP_6680_elements(526);
    -- CP-element group 528:  transition  input  no-bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	527 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	531 
    -- CP-element group 528:  members (2) 
      -- CP-element group 528: 	 branch_block_stmt_1353/if_stmt_2054_if_link/$exit
      -- CP-element group 528: 	 branch_block_stmt_1353/if_stmt_2054_if_link/if_choice_transition
      -- 
    if_choice_transition_9665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2054_branch_ack_1, ack => minSumDecode_CP_6680_elements(528)); -- 
    -- CP-element group 529:  transition  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	526 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	530 
    -- CP-element group 529:  members (1) 
      -- CP-element group 529: 	 branch_block_stmt_1353/if_stmt_2054_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(529) <= minSumDecode_CP_6680_elements(526);
    -- CP-element group 530:  transition  input  no-bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	529 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (2) 
      -- CP-element group 530: 	 branch_block_stmt_1353/if_stmt_2054_else_link/$exit
      -- CP-element group 530: 	 branch_block_stmt_1353/if_stmt_2054_else_link/else_choice_transition
      -- 
    else_choice_transition_9669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2054_branch_ack_0, ack => minSumDecode_CP_6680_elements(530)); -- 
    -- CP-element group 531:  place  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	528 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	1022 
    -- CP-element group 531:  members (1) 
      -- CP-element group 531: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread
      -- 
    minSumDecode_CP_6680_elements(531) <= minSumDecode_CP_6680_elements(528);
    -- CP-element group 532:  place  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	1029 
    -- CP-element group 532:  members (1) 
      -- CP-element group 532: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_bbx_xnphx_xi43
      -- 
    minSumDecode_CP_6680_elements(532) <= minSumDecode_CP_6680_elements(530);
    -- CP-element group 533:  fork  transition  output  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	51 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533: 	535 
    -- CP-element group 533:  members (17) 
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/STORE_Nitr_required_2066_Split/split_ack
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_root_address_calculated
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_word_address_calculated
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/STORE_Nitr_required_2066_Split/split_req
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_update_start_
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_sample_start_
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/STORE_Nitr_required_2066_Split/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/STORE_Nitr_required_2066_Split/$exit
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/word_0/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/word_0/rr
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/word_0/$entry
      -- CP-element group 533: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/word_0/cr
      -- 
    cr_9706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(533), ack => STORE_Nitr_required_2066_store_0_req_1); -- 
    rr_9695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(533), ack => STORE_Nitr_required_2066_store_0_req_0); -- 
    minSumDecode_CP_6680_elements(533) <= minSumDecode_CP_6680_elements(51);
    -- CP-element group 534:  transition  input  no-bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534:  members (5) 
      -- CP-element group 534: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/$exit
      -- CP-element group 534: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_sample_completed_
      -- CP-element group 534: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/$exit
      -- CP-element group 534: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/word_0/$exit
      -- CP-element group 534: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Sample/word_access_start/word_0/ra
      -- 
    ra_9696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_Nitr_required_2066_store_0_ack_0, ack => minSumDecode_CP_6680_elements(534)); -- 
    -- CP-element group 535:  transition  input  no-bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	533 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	52 
    -- CP-element group 535:  members (6) 
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_update_completed_
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/$exit
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/$exit
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/$exit
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/word_0/$exit
      -- CP-element group 535: 	 branch_block_stmt_1353/assign_stmt_2068/STORE_Nitr_required_2066_Update/word_access_complete/word_0/ca
      -- 
    ca_9707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_Nitr_required_2066_store_0_ack_1, ack => minSumDecode_CP_6680_elements(535)); -- 
    -- CP-element group 536:  fork  transition  output  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	53 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	537 
    -- CP-element group 536: 	538 
    -- CP-element group 536: 	539 
    -- CP-element group 536: 	540 
    -- CP-element group 536: 	542 
    -- CP-element group 536: 	544 
    -- CP-element group 536: 	547 
    -- CP-element group 536:  members (22) 
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Sample/rr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Sample/rr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_complete/req
      -- 
    rr_9718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => UGT_u16_u1_2075_inst_req_0); -- 
    cr_9723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => UGT_u16_u1_2075_inst_req_1); -- 
    rr_9732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => ADD_u16_u16_2081_inst_req_0); -- 
    cr_9737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => ADD_u16_u16_2081_inst_req_1); -- 
    cr_9751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => type_cast_2085_inst_req_1); -- 
    cr_9765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => ADD_u64_u64_2091_inst_req_1); -- 
    req_9779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(536), ack => MUX_2098_inst_req_1); -- 
    minSumDecode_CP_6680_elements(536) <= minSumDecode_CP_6680_elements(53);
    -- CP-element group 537:  transition  input  no-bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	536 
    -- CP-element group 537: successors 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_sample_completed_
      -- CP-element group 537: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Sample/$exit
      -- CP-element group 537: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Sample/ra
      -- 
    ra_9719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_2075_inst_ack_0, ack => minSumDecode_CP_6680_elements(537)); -- 
    -- CP-element group 538:  transition  input  no-bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	536 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	545 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_update_completed_
      -- CP-element group 538: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Update/$exit
      -- CP-element group 538: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/UGT_u16_u1_2075_Update/ca
      -- 
    ca_9724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_2075_inst_ack_1, ack => minSumDecode_CP_6680_elements(538)); -- 
    -- CP-element group 539:  transition  input  no-bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	536 
    -- CP-element group 539: successors 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Sample/ra
      -- 
    ra_9733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2081_inst_ack_0, ack => minSumDecode_CP_6680_elements(539)); -- 
    -- CP-element group 540:  transition  input  output  no-bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	536 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540:  members (6) 
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u16_u16_2081_Update/ca
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_sample_start_
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Sample/$entry
      -- CP-element group 540: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Sample/rr
      -- 
    ca_9738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2081_inst_ack_1, ack => minSumDecode_CP_6680_elements(540)); -- 
    rr_9746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(540), ack => type_cast_2085_inst_req_0); -- 
    -- CP-element group 541:  transition  input  no-bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	540 
    -- CP-element group 541: successors 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_sample_completed_
      -- CP-element group 541: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Sample/$exit
      -- CP-element group 541: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Sample/ra
      -- 
    ra_9747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2085_inst_ack_0, ack => minSumDecode_CP_6680_elements(541)); -- 
    -- CP-element group 542:  transition  input  output  no-bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	536 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542:  members (6) 
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_update_completed_
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Update/$exit
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/type_cast_2085_Update/ca
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_sample_start_
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Sample/$entry
      -- CP-element group 542: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Sample/rr
      -- 
    ca_9752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2085_inst_ack_1, ack => minSumDecode_CP_6680_elements(542)); -- 
    rr_9760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(542), ack => ADD_u64_u64_2091_inst_req_0); -- 
    -- CP-element group 543:  transition  input  no-bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	542 
    -- CP-element group 543: successors 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_sample_completed_
      -- CP-element group 543: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Sample/$exit
      -- CP-element group 543: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Sample/ra
      -- 
    ra_9761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2091_inst_ack_0, ack => minSumDecode_CP_6680_elements(543)); -- 
    -- CP-element group 544:  transition  input  no-bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	536 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	545 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_update_completed_
      -- CP-element group 544: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Update/$exit
      -- CP-element group 544: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/ADD_u64_u64_2091_Update/ca
      -- 
    ca_9766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2091_inst_ack_1, ack => minSumDecode_CP_6680_elements(544)); -- 
    -- CP-element group 545:  join  transition  output  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	538 
    -- CP-element group 545: 	544 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	546 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_sample_start_
      -- CP-element group 545: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_start/$entry
      -- CP-element group 545: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_start/req
      -- 
    req_9774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(545), ack => MUX_2098_inst_req_0); -- 
    minSumDecode_cp_element_group_545: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_545"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(538) & minSumDecode_CP_6680_elements(544);
      gj_minSumDecode_cp_element_group_545 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(545), clk => clk, reset => reset); --
    end block;
    -- CP-element group 546:  transition  input  no-bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	545 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	548 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_sample_completed_
      -- CP-element group 546: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_start/$exit
      -- CP-element group 546: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_start/ack
      -- 
    ack_9775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2098_inst_ack_0, ack => minSumDecode_CP_6680_elements(546)); -- 
    -- CP-element group 547:  transition  input  no-bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	536 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	548 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_update_completed_
      -- CP-element group 547: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_complete/$exit
      -- CP-element group 547: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/MUX_2098_complete/ack
      -- 
    ack_9780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2098_inst_ack_1, ack => minSumDecode_CP_6680_elements(547)); -- 
    -- CP-element group 548:  join  transition  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	546 
    -- CP-element group 548: 	547 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	54 
    -- CP-element group 548:  members (1) 
      -- CP-element group 548: 	 branch_block_stmt_1353/assign_stmt_2076_to_assign_stmt_2099/$exit
      -- 
    minSumDecode_cp_element_group_548: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_548"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(546) & minSumDecode_CP_6680_elements(547);
      gj_minSumDecode_cp_element_group_548 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(548), clk => clk, reset => reset); --
    end block;
    -- CP-element group 549:  fork  transition  output  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	55 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	550 
    -- CP-element group 549: 	551 
    -- CP-element group 549: 	552 
    -- CP-element group 549: 	553 
    -- CP-element group 549: 	555 
    -- CP-element group 549: 	557 
    -- CP-element group 549: 	559 
    -- CP-element group 549:  members (66) 
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_sample_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_update_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_root_address_calculated
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_offset_calculated
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_resized_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_scaled_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_computed_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_resize_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_resize_0/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_resize_0/index_resize_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_resize_0/index_resize_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_scale_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_scale_0/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_scale_0/scale_rename_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_index_scale_0/scale_rename_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_final_index_sum_regn/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_final_index_sum_regn/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_final_index_sum_regn/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_final_index_sum_regn/ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_base_plus_offset/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_base_plus_offset/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_base_plus_offset/sum_rename_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2119_base_plus_offset/sum_rename_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_request/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_request/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_complete/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_complete/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_sample_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_update_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_root_address_calculated
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_offset_calculated
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_resized_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_scaled_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_computed_0
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_resize_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_resize_0/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_resize_0/index_resize_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_resize_0/index_resize_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_scale_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_scale_0/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_scale_0/scale_rename_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_index_scale_0/scale_rename_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_final_index_sum_regn/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_final_index_sum_regn/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_final_index_sum_regn/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_final_index_sum_regn/ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_base_plus_offset/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_base_plus_offset/$exit
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_base_plus_offset/sum_rename_req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/array_obj_ref_2124_base_plus_offset/sum_rename_ack
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_request/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_request/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_complete/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_complete/req
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_update_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/word_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/word_0/cr
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_update_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Update/cr
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_update_start_
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Update/cr
      -- 
    req_9821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => addr_of_2120_final_reg_req_1); -- 
    req_9816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => addr_of_2120_final_reg_req_0); -- 
    req_9860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => addr_of_2125_final_reg_req_1); -- 
    req_9855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => addr_of_2125_final_reg_req_0); -- 
    cr_9905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => ptr_deref_2129_load_0_req_1); -- 
    cr_9924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => type_cast_2133_inst_req_1); -- 
    cr_9938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(549), ack => SGT_f64_u1_2139_inst_req_1); -- 
    minSumDecode_CP_6680_elements(549) <= minSumDecode_CP_6680_elements(55);
    -- CP-element group 550:  transition  input  no-bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	549 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	560 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_sample_completed_
      -- CP-element group 550: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_request/$exit
      -- CP-element group 550: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_request/ack
      -- 
    ack_9817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2120_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(550)); -- 
    -- CP-element group 551:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	549 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	554 
    -- CP-element group 551:  members (24) 
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_update_completed_
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_complete/$exit
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2120_complete/ack
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_sample_start_
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_address_calculated
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_word_address_calculated
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_root_address_calculated
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_address_resized
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_addr_resize/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_addr_resize/$exit
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_addr_resize/base_resize_req
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_addr_resize/base_resize_ack
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_plus_offset/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_plus_offset/$exit
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_plus_offset/sum_rename_req
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_base_plus_offset/sum_rename_ack
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_word_addrgen/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_word_addrgen/$exit
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_word_addrgen/root_register_req
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_word_addrgen/root_register_ack
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/word_0/$entry
      -- CP-element group 551: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/word_0/rr
      -- 
    ack_9822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 551_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2120_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(551)); -- 
    rr_9894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(551), ack => ptr_deref_2129_load_0_req_0); -- 
    -- CP-element group 552:  transition  input  no-bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	549 
    -- CP-element group 552: successors 
    -- CP-element group 552: 	560 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_request/$exit
      -- CP-element group 552: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_request/ack
      -- 
    ack_9856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2125_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(552)); -- 
    -- CP-element group 553:  transition  input  no-bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	549 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	560 
    -- CP-element group 553:  members (3) 
      -- CP-element group 553: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_complete/$exit
      -- CP-element group 553: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/addr_of_2125_complete/ack
      -- 
    ack_9861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2125_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(553)); -- 
    -- CP-element group 554:  transition  input  no-bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	551 
    -- CP-element group 554: successors 
    -- CP-element group 554:  members (5) 
      -- CP-element group 554: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_sample_completed_
      -- CP-element group 554: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/$exit
      -- CP-element group 554: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/$exit
      -- CP-element group 554: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/word_0/$exit
      -- CP-element group 554: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Sample/word_access_start/word_0/ra
      -- 
    ra_9895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2129_load_0_ack_0, ack => minSumDecode_CP_6680_elements(554)); -- 
    -- CP-element group 555:  transition  input  output  no-bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	549 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	556 
    -- CP-element group 555:  members (12) 
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_update_completed_
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/$exit
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/$exit
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/word_0/$exit
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/word_access_complete/word_0/ca
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/ptr_deref_2129_Merge/$entry
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/ptr_deref_2129_Merge/$exit
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/ptr_deref_2129_Merge/merge_req
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/ptr_deref_2129_Update/ptr_deref_2129_Merge/merge_ack
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_sample_start_
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Sample/$entry
      -- CP-element group 555: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Sample/rr
      -- 
    ca_9906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2129_load_0_ack_1, ack => minSumDecode_CP_6680_elements(555)); -- 
    rr_9919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(555), ack => type_cast_2133_inst_req_0); -- 
    -- CP-element group 556:  transition  input  no-bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	555 
    -- CP-element group 556: successors 
    -- CP-element group 556:  members (3) 
      -- CP-element group 556: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_sample_completed_
      -- CP-element group 556: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Sample/ra
      -- 
    ra_9920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_0, ack => minSumDecode_CP_6680_elements(556)); -- 
    -- CP-element group 557:  transition  input  output  no-bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	549 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557:  members (6) 
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_update_completed_
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/type_cast_2133_Update/ca
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_sample_start_
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Sample/$entry
      -- CP-element group 557: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Sample/rr
      -- 
    ca_9925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_1, ack => minSumDecode_CP_6680_elements(557)); -- 
    rr_9933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(557), ack => SGT_f64_u1_2139_inst_req_0); -- 
    -- CP-element group 558:  transition  input  no-bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	557 
    -- CP-element group 558: successors 
    -- CP-element group 558:  members (3) 
      -- CP-element group 558: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_sample_completed_
      -- CP-element group 558: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Sample/$exit
      -- CP-element group 558: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Sample/ra
      -- 
    ra_9934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 558_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2139_inst_ack_0, ack => minSumDecode_CP_6680_elements(558)); -- 
    -- CP-element group 559:  transition  input  no-bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	549 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	560 
    -- CP-element group 559:  members (3) 
      -- CP-element group 559: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_update_completed_
      -- CP-element group 559: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Update/$exit
      -- CP-element group 559: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/SGT_f64_u1_2139_Update/ca
      -- 
    ca_9939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2139_inst_ack_1, ack => minSumDecode_CP_6680_elements(559)); -- 
    -- CP-element group 560:  join  transition  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	550 
    -- CP-element group 560: 	552 
    -- CP-element group 560: 	553 
    -- CP-element group 560: 	559 
    -- CP-element group 560: successors 
    -- CP-element group 560: 	56 
    -- CP-element group 560:  members (1) 
      -- CP-element group 560: 	 branch_block_stmt_1353/assign_stmt_2121_to_assign_stmt_2140/$exit
      -- 
    minSumDecode_cp_element_group_560: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_560"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(550) & minSumDecode_CP_6680_elements(552) & minSumDecode_CP_6680_elements(553) & minSumDecode_CP_6680_elements(559);
      gj_minSumDecode_cp_element_group_560 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(560), clk => clk, reset => reset); --
    end block;
    -- CP-element group 561:  transition  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	56 
    -- CP-element group 561: successors 
    -- CP-element group 561:  members (1) 
      -- CP-element group 561: 	 branch_block_stmt_1353/if_stmt_2141_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(561) <= minSumDecode_CP_6680_elements(56);
    -- CP-element group 562:  transition  output  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	56 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	563 
    -- CP-element group 562:  members (3) 
      -- CP-element group 562: 	 branch_block_stmt_1353/if_stmt_2141_eval_test/$entry
      -- CP-element group 562: 	 branch_block_stmt_1353/if_stmt_2141_eval_test/$exit
      -- CP-element group 562: 	 branch_block_stmt_1353/if_stmt_2141_eval_test/branch_req
      -- 
    branch_req_9947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(562), ack => if_stmt_2141_branch_req_0); -- 
    minSumDecode_CP_6680_elements(562) <= minSumDecode_CP_6680_elements(56);
    -- CP-element group 563:  branch  place  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	562 
    -- CP-element group 563: successors 
    -- CP-element group 563: 	564 
    -- CP-element group 563: 	566 
    -- CP-element group 563:  members (1) 
      -- CP-element group 563: 	 branch_block_stmt_1353/R_iNsTr_108_2142_place
      -- 
    minSumDecode_CP_6680_elements(563) <= minSumDecode_CP_6680_elements(562);
    -- CP-element group 564:  transition  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	563 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	565 
    -- CP-element group 564:  members (1) 
      -- CP-element group 564: 	 branch_block_stmt_1353/if_stmt_2141_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(564) <= minSumDecode_CP_6680_elements(563);
    -- CP-element group 565:  transition  input  no-bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	564 
    -- CP-element group 565: successors 
    -- CP-element group 565: 	568 
    -- CP-element group 565:  members (2) 
      -- CP-element group 565: 	 branch_block_stmt_1353/if_stmt_2141_if_link/$exit
      -- CP-element group 565: 	 branch_block_stmt_1353/if_stmt_2141_if_link/if_choice_transition
      -- 
    if_choice_transition_9952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2141_branch_ack_1, ack => minSumDecode_CP_6680_elements(565)); -- 
    -- CP-element group 566:  transition  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	563 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	567 
    -- CP-element group 566:  members (1) 
      -- CP-element group 566: 	 branch_block_stmt_1353/if_stmt_2141_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(566) <= minSumDecode_CP_6680_elements(563);
    -- CP-element group 567:  transition  input  no-bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	566 
    -- CP-element group 567: successors 
    -- CP-element group 567: 	569 
    -- CP-element group 567:  members (2) 
      -- CP-element group 567: 	 branch_block_stmt_1353/if_stmt_2141_else_link/$exit
      -- CP-element group 567: 	 branch_block_stmt_1353/if_stmt_2141_else_link/else_choice_transition
      -- 
    else_choice_transition_9956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2141_branch_ack_0, ack => minSumDecode_CP_6680_elements(567)); -- 
    -- CP-element group 568:  place  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	565 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	1051 
    -- CP-element group 568:  members (1) 
      -- CP-element group 568: 	 branch_block_stmt_1353/bb_29_bb_30
      -- 
    minSumDecode_CP_6680_elements(568) <= minSumDecode_CP_6680_elements(565);
    -- CP-element group 569:  place  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	567 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	1067 
    -- CP-element group 569:  members (1) 
      -- CP-element group 569: 	 branch_block_stmt_1353/bb_29_bb_33
      -- 
    minSumDecode_CP_6680_elements(569) <= minSumDecode_CP_6680_elements(567);
    -- CP-element group 570:  join  fork  transition  output  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	57 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	571 
    -- CP-element group 570: 	572 
    -- CP-element group 570: 	574 
    -- CP-element group 570: 	576 
    -- CP-element group 570:  members (33) 
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_sample_start_
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_update_start_
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_address_calculated
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_word_address_calculated
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_root_address_calculated
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_address_resized
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_addr_resize/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_addr_resize/$exit
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_addr_resize/base_resize_req
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_addr_resize/base_resize_ack
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_plus_offset/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_plus_offset/$exit
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_plus_offset/sum_rename_req
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_base_plus_offset/sum_rename_ack
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_word_addrgen/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_word_addrgen/$exit
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_word_addrgen/root_register_req
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_word_addrgen/root_register_ack
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/word_0/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/word_0/rr
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/word_0/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/word_0/cr
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_update_start_
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Update/cr
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_update_start_
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Update/cr
      -- 
    cr_10005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(570), ack => ptr_deref_2150_load_0_req_1); -- 
    rr_9994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(570), ack => ptr_deref_2150_load_0_req_0); -- 
    cr_10024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(570), ack => type_cast_2154_inst_req_1); -- 
    cr_10038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(570), ack => SGT_f64_u1_2160_inst_req_1); -- 
    minSumDecode_CP_6680_elements(570) <= minSumDecode_CP_6680_elements(57);
    -- CP-element group 571:  transition  input  no-bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	570 
    -- CP-element group 571: successors 
    -- CP-element group 571:  members (5) 
      -- CP-element group 571: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/$exit
      -- CP-element group 571: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/$exit
      -- CP-element group 571: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/word_0/$exit
      -- CP-element group 571: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Sample/word_access_start/word_0/ra
      -- 
    ra_9995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2150_load_0_ack_0, ack => minSumDecode_CP_6680_elements(571)); -- 
    -- CP-element group 572:  transition  input  output  no-bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	570 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	573 
    -- CP-element group 572:  members (12) 
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/$exit
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/$exit
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/word_0/$exit
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/word_access_complete/word_0/ca
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/ptr_deref_2150_Merge/$entry
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/ptr_deref_2150_Merge/$exit
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/ptr_deref_2150_Merge/merge_req
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/ptr_deref_2150_Update/ptr_deref_2150_Merge/merge_ack
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_sample_start_
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Sample/$entry
      -- CP-element group 572: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Sample/rr
      -- 
    ca_10006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2150_load_0_ack_1, ack => minSumDecode_CP_6680_elements(572)); -- 
    rr_10019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(572), ack => type_cast_2154_inst_req_0); -- 
    -- CP-element group 573:  transition  input  no-bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	572 
    -- CP-element group 573: successors 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_sample_completed_
      -- CP-element group 573: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Sample/$exit
      -- CP-element group 573: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Sample/ra
      -- 
    ra_10020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2154_inst_ack_0, ack => minSumDecode_CP_6680_elements(573)); -- 
    -- CP-element group 574:  transition  input  output  no-bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	570 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	575 
    -- CP-element group 574:  members (6) 
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_update_completed_
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Update/$exit
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/type_cast_2154_Update/ca
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_sample_start_
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Sample/$entry
      -- CP-element group 574: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Sample/rr
      -- 
    ca_10025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2154_inst_ack_1, ack => minSumDecode_CP_6680_elements(574)); -- 
    rr_10033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(574), ack => SGT_f64_u1_2160_inst_req_0); -- 
    -- CP-element group 575:  transition  input  no-bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	574 
    -- CP-element group 575: successors 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_sample_completed_
      -- CP-element group 575: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Sample/$exit
      -- CP-element group 575: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Sample/ra
      -- 
    ra_10034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2160_inst_ack_0, ack => minSumDecode_CP_6680_elements(575)); -- 
    -- CP-element group 576:  transition  input  no-bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	570 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	58 
    -- CP-element group 576:  members (4) 
      -- CP-element group 576: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/$exit
      -- CP-element group 576: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_update_completed_
      -- CP-element group 576: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Update/$exit
      -- CP-element group 576: 	 branch_block_stmt_1353/assign_stmt_2151_to_assign_stmt_2161/SGT_f64_u1_2160_Update/ca
      -- 
    ca_10039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SGT_f64_u1_2160_inst_ack_1, ack => minSumDecode_CP_6680_elements(576)); -- 
    -- CP-element group 577:  transition  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	58 
    -- CP-element group 577: successors 
    -- CP-element group 577:  members (1) 
      -- CP-element group 577: 	 branch_block_stmt_1353/if_stmt_2162_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(577) <= minSumDecode_CP_6680_elements(58);
    -- CP-element group 578:  transition  output  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	58 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	579 
    -- CP-element group 578:  members (3) 
      -- CP-element group 578: 	 branch_block_stmt_1353/if_stmt_2162_eval_test/$entry
      -- CP-element group 578: 	 branch_block_stmt_1353/if_stmt_2162_eval_test/$exit
      -- CP-element group 578: 	 branch_block_stmt_1353/if_stmt_2162_eval_test/branch_req
      -- 
    branch_req_10047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(578), ack => if_stmt_2162_branch_req_0); -- 
    minSumDecode_CP_6680_elements(578) <= minSumDecode_CP_6680_elements(58);
    -- CP-element group 579:  branch  place  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	578 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	580 
    -- CP-element group 579: 	582 
    -- CP-element group 579:  members (1) 
      -- CP-element group 579: 	 branch_block_stmt_1353/R_iNsTr_113_2163_place
      -- 
    minSumDecode_CP_6680_elements(579) <= minSumDecode_CP_6680_elements(578);
    -- CP-element group 580:  transition  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	579 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	581 
    -- CP-element group 580:  members (1) 
      -- CP-element group 580: 	 branch_block_stmt_1353/if_stmt_2162_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(580) <= minSumDecode_CP_6680_elements(579);
    -- CP-element group 581:  transition  input  no-bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	580 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	584 
    -- CP-element group 581:  members (2) 
      -- CP-element group 581: 	 branch_block_stmt_1353/if_stmt_2162_if_link/$exit
      -- CP-element group 581: 	 branch_block_stmt_1353/if_stmt_2162_if_link/if_choice_transition
      -- 
    if_choice_transition_10052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 581_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2162_branch_ack_1, ack => minSumDecode_CP_6680_elements(581)); -- 
    -- CP-element group 582:  transition  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	579 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	583 
    -- CP-element group 582:  members (1) 
      -- CP-element group 582: 	 branch_block_stmt_1353/if_stmt_2162_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(582) <= minSumDecode_CP_6680_elements(579);
    -- CP-element group 583:  transition  input  no-bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	582 
    -- CP-element group 583: successors 
    -- CP-element group 583: 	585 
    -- CP-element group 583:  members (2) 
      -- CP-element group 583: 	 branch_block_stmt_1353/if_stmt_2162_else_link/$exit
      -- CP-element group 583: 	 branch_block_stmt_1353/if_stmt_2162_else_link/else_choice_transition
      -- 
    else_choice_transition_10056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2162_branch_ack_0, ack => minSumDecode_CP_6680_elements(583)); -- 
    -- CP-element group 584:  place  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	581 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	1054 
    -- CP-element group 584:  members (1) 
      -- CP-element group 584: 	 branch_block_stmt_1353/bb_30_bb_31
      -- 
    minSumDecode_CP_6680_elements(584) <= minSumDecode_CP_6680_elements(581);
    -- CP-element group 585:  place  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	583 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	1057 
    -- CP-element group 585:  members (1) 
      -- CP-element group 585: 	 branch_block_stmt_1353/bb_30_bb_32
      -- 
    minSumDecode_CP_6680_elements(585) <= minSumDecode_CP_6680_elements(583);
    -- CP-element group 586:  fork  transition  output  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	59 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	587 
    -- CP-element group 586: 	588 
    -- CP-element group 586:  members (17) 
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_sample_start_
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_update_start_
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_word_address_calculated
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_root_address_calculated
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/STORE_is_decoded_2169_Split/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/STORE_is_decoded_2169_Split/$exit
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/STORE_is_decoded_2169_Split/split_req
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/STORE_is_decoded_2169_Split/split_ack
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/word_0/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/word_0/rr
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/word_0/$entry
      -- CP-element group 586: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/word_0/cr
      -- 
    cr_10093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(586), ack => STORE_is_decoded_2169_store_0_req_1); -- 
    rr_10082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(586), ack => STORE_is_decoded_2169_store_0_req_0); -- 
    minSumDecode_CP_6680_elements(586) <= minSumDecode_CP_6680_elements(59);
    -- CP-element group 587:  transition  input  no-bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	586 
    -- CP-element group 587: successors 
    -- CP-element group 587:  members (5) 
      -- CP-element group 587: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_sample_completed_
      -- CP-element group 587: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/$exit
      -- CP-element group 587: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/$exit
      -- CP-element group 587: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/word_0/$exit
      -- CP-element group 587: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Sample/word_access_start/word_0/ra
      -- 
    ra_10083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 587_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2169_store_0_ack_0, ack => minSumDecode_CP_6680_elements(587)); -- 
    -- CP-element group 588:  transition  input  no-bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	586 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	60 
    -- CP-element group 588:  members (6) 
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/$exit
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_update_completed_
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/$exit
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/$exit
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/word_0/$exit
      -- CP-element group 588: 	 branch_block_stmt_1353/assign_stmt_2172/STORE_is_decoded_2169_Update/word_access_complete/word_0/ca
      -- 
    ca_10094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2169_store_0_ack_1, ack => minSumDecode_CP_6680_elements(588)); -- 
    -- CP-element group 589:  join  fork  transition  output  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	61 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	590 
    -- CP-element group 589: 	591 
    -- CP-element group 589:  members (31) 
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_sample_start_
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_update_start_
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_address_calculated
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_word_address_calculated
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_root_address_calculated
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_address_resized
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_addr_resize/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_addr_resize/$exit
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_addr_resize/base_resize_req
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_addr_resize/base_resize_ack
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_plus_offset/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_plus_offset/$exit
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_plus_offset/sum_rename_req
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_base_plus_offset/sum_rename_ack
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_word_addrgen/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_word_addrgen/$exit
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_word_addrgen/root_register_req
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_word_addrgen/root_register_ack
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/ptr_deref_2184_Split/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/ptr_deref_2184_Split/$exit
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/ptr_deref_2184_Split/split_req
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/ptr_deref_2184_Split/split_ack
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/word_0/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/word_0/rr
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/word_0/$entry
      -- CP-element group 589: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/word_0/cr
      -- 
    cr_10146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(589), ack => ptr_deref_2184_store_0_req_1); -- 
    rr_10135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(589), ack => ptr_deref_2184_store_0_req_0); -- 
    minSumDecode_CP_6680_elements(589) <= minSumDecode_CP_6680_elements(61);
    -- CP-element group 590:  transition  input  no-bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	589 
    -- CP-element group 590: successors 
    -- CP-element group 590:  members (5) 
      -- CP-element group 590: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_sample_completed_
      -- CP-element group 590: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/$exit
      -- CP-element group 590: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/$exit
      -- CP-element group 590: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/word_0/$exit
      -- CP-element group 590: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Sample/word_access_start/word_0/ra
      -- 
    ra_10136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 590_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2184_store_0_ack_0, ack => minSumDecode_CP_6680_elements(590)); -- 
    -- CP-element group 591:  transition  input  no-bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	589 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	62 
    -- CP-element group 591:  members (6) 
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/$exit
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_update_completed_
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/$exit
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/$exit
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/word_0/$exit
      -- CP-element group 591: 	 branch_block_stmt_1353/assign_stmt_2187/ptr_deref_2184_Update/word_access_complete/word_0/ca
      -- 
    ca_10147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2184_store_0_ack_1, ack => minSumDecode_CP_6680_elements(591)); -- 
    -- CP-element group 592:  fork  transition  output  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	63 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	593 
    -- CP-element group 592: 	594 
    -- CP-element group 592:  members (7) 
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/$entry
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_sample_start_
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_update_start_
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Sample/$entry
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Sample/rr
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Update/$entry
      -- CP-element group 592: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Update/cr
      -- 
    rr_10158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(592), ack => SLT_f64_u1_2194_inst_req_0); -- 
    cr_10163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(592), ack => SLT_f64_u1_2194_inst_req_1); -- 
    minSumDecode_CP_6680_elements(592) <= minSumDecode_CP_6680_elements(63);
    -- CP-element group 593:  transition  input  no-bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	592 
    -- CP-element group 593: successors 
    -- CP-element group 593:  members (3) 
      -- CP-element group 593: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_sample_completed_
      -- CP-element group 593: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Sample/$exit
      -- CP-element group 593: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Sample/ra
      -- 
    ra_10159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 593_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2194_inst_ack_0, ack => minSumDecode_CP_6680_elements(593)); -- 
    -- CP-element group 594:  transition  input  no-bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	592 
    -- CP-element group 594: successors 
    -- CP-element group 594: 	64 
    -- CP-element group 594:  members (4) 
      -- CP-element group 594: 	 branch_block_stmt_1353/assign_stmt_2195/$exit
      -- CP-element group 594: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_update_completed_
      -- CP-element group 594: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Update/$exit
      -- CP-element group 594: 	 branch_block_stmt_1353/assign_stmt_2195/SLT_f64_u1_2194_Update/ca
      -- 
    ca_10164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 594_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2194_inst_ack_1, ack => minSumDecode_CP_6680_elements(594)); -- 
    -- CP-element group 595:  transition  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	64 
    -- CP-element group 595: successors 
    -- CP-element group 595:  members (1) 
      -- CP-element group 595: 	 branch_block_stmt_1353/if_stmt_2196_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(595) <= minSumDecode_CP_6680_elements(64);
    -- CP-element group 596:  transition  output  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	64 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	597 
    -- CP-element group 596:  members (3) 
      -- CP-element group 596: 	 branch_block_stmt_1353/if_stmt_2196_eval_test/$entry
      -- CP-element group 596: 	 branch_block_stmt_1353/if_stmt_2196_eval_test/$exit
      -- CP-element group 596: 	 branch_block_stmt_1353/if_stmt_2196_eval_test/branch_req
      -- 
    branch_req_10172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(596), ack => if_stmt_2196_branch_req_0); -- 
    minSumDecode_CP_6680_elements(596) <= minSumDecode_CP_6680_elements(64);
    -- CP-element group 597:  branch  place  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	596 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	598 
    -- CP-element group 597: 	600 
    -- CP-element group 597:  members (1) 
      -- CP-element group 597: 	 branch_block_stmt_1353/R_iNsTr_115_2197_place
      -- 
    minSumDecode_CP_6680_elements(597) <= minSumDecode_CP_6680_elements(596);
    -- CP-element group 598:  transition  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	597 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	599 
    -- CP-element group 598:  members (1) 
      -- CP-element group 598: 	 branch_block_stmt_1353/if_stmt_2196_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(598) <= minSumDecode_CP_6680_elements(597);
    -- CP-element group 599:  transition  input  no-bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	598 
    -- CP-element group 599: successors 
    -- CP-element group 599: 	602 
    -- CP-element group 599:  members (2) 
      -- CP-element group 599: 	 branch_block_stmt_1353/if_stmt_2196_if_link/$exit
      -- CP-element group 599: 	 branch_block_stmt_1353/if_stmt_2196_if_link/if_choice_transition
      -- 
    if_choice_transition_10177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 599_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2196_branch_ack_1, ack => minSumDecode_CP_6680_elements(599)); -- 
    -- CP-element group 600:  transition  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	597 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	601 
    -- CP-element group 600:  members (1) 
      -- CP-element group 600: 	 branch_block_stmt_1353/if_stmt_2196_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(600) <= minSumDecode_CP_6680_elements(597);
    -- CP-element group 601:  transition  input  no-bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	600 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (2) 
      -- CP-element group 601: 	 branch_block_stmt_1353/if_stmt_2196_else_link/$exit
      -- CP-element group 601: 	 branch_block_stmt_1353/if_stmt_2196_else_link/else_choice_transition
      -- 
    else_choice_transition_10181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2196_branch_ack_0, ack => minSumDecode_CP_6680_elements(601)); -- 
    -- CP-element group 602:  place  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	599 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	1070 
    -- CP-element group 602:  members (1) 
      -- CP-element group 602: 	 branch_block_stmt_1353/bb_33_bb_34
      -- 
    minSumDecode_CP_6680_elements(602) <= minSumDecode_CP_6680_elements(599);
    -- CP-element group 603:  place  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	601 
    -- CP-element group 603: successors 
    -- CP-element group 603: 	1090 
    -- CP-element group 603:  members (1) 
      -- CP-element group 603: 	 branch_block_stmt_1353/bb_33_bb_37
      -- 
    minSumDecode_CP_6680_elements(603) <= minSumDecode_CP_6680_elements(601);
    -- CP-element group 604:  join  fork  transition  output  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	65 
    -- CP-element group 604: successors 
    -- CP-element group 604: 	605 
    -- CP-element group 604: 	606 
    -- CP-element group 604: 	608 
    -- CP-element group 604: 	610 
    -- CP-element group 604:  members (33) 
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_sample_start_
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_update_start_
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_address_calculated
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_word_address_calculated
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_root_address_calculated
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_address_resized
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_addr_resize/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_addr_resize/$exit
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_addr_resize/base_resize_req
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_addr_resize/base_resize_ack
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_plus_offset/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_plus_offset/$exit
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_plus_offset/sum_rename_req
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_base_plus_offset/sum_rename_ack
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_word_addrgen/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_word_addrgen/$exit
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_word_addrgen/root_register_req
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_word_addrgen/root_register_ack
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/word_0/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/word_0/rr
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/word_0/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/word_0/cr
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_update_start_
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Update/cr
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_update_start_
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Update/cr
      -- 
    cr_10230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(604), ack => ptr_deref_2205_load_0_req_1); -- 
    rr_10219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(604), ack => ptr_deref_2205_load_0_req_0); -- 
    cr_10249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(604), ack => type_cast_2209_inst_req_1); -- 
    cr_10263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(604), ack => SLT_f64_u1_2215_inst_req_1); -- 
    minSumDecode_CP_6680_elements(604) <= minSumDecode_CP_6680_elements(65);
    -- CP-element group 605:  transition  input  no-bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	604 
    -- CP-element group 605: successors 
    -- CP-element group 605:  members (5) 
      -- CP-element group 605: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_sample_completed_
      -- CP-element group 605: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/$exit
      -- CP-element group 605: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/$exit
      -- CP-element group 605: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/word_0/$exit
      -- CP-element group 605: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Sample/word_access_start/word_0/ra
      -- 
    ra_10220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 605_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2205_load_0_ack_0, ack => minSumDecode_CP_6680_elements(605)); -- 
    -- CP-element group 606:  transition  input  output  no-bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	604 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	607 
    -- CP-element group 606:  members (12) 
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_update_completed_
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/$exit
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/$exit
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/word_0/$exit
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/word_access_complete/word_0/ca
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/ptr_deref_2205_Merge/$entry
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/ptr_deref_2205_Merge/$exit
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/ptr_deref_2205_Merge/merge_req
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/ptr_deref_2205_Update/ptr_deref_2205_Merge/merge_ack
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_sample_start_
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Sample/$entry
      -- CP-element group 606: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Sample/rr
      -- 
    ca_10231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2205_load_0_ack_1, ack => minSumDecode_CP_6680_elements(606)); -- 
    rr_10244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(606), ack => type_cast_2209_inst_req_0); -- 
    -- CP-element group 607:  transition  input  no-bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	606 
    -- CP-element group 607: successors 
    -- CP-element group 607:  members (3) 
      -- CP-element group 607: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_sample_completed_
      -- CP-element group 607: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Sample/$exit
      -- CP-element group 607: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Sample/ra
      -- 
    ra_10245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2209_inst_ack_0, ack => minSumDecode_CP_6680_elements(607)); -- 
    -- CP-element group 608:  transition  input  output  no-bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	604 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	609 
    -- CP-element group 608:  members (6) 
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_update_completed_
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Update/$exit
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/type_cast_2209_Update/ca
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_sample_start_
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Sample/$entry
      -- CP-element group 608: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Sample/rr
      -- 
    ca_10250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2209_inst_ack_1, ack => minSumDecode_CP_6680_elements(608)); -- 
    rr_10258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(608), ack => SLT_f64_u1_2215_inst_req_0); -- 
    -- CP-element group 609:  transition  input  no-bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	608 
    -- CP-element group 609: successors 
    -- CP-element group 609:  members (3) 
      -- CP-element group 609: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_sample_completed_
      -- CP-element group 609: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Sample/$exit
      -- CP-element group 609: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Sample/ra
      -- 
    ra_10259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2215_inst_ack_0, ack => minSumDecode_CP_6680_elements(609)); -- 
    -- CP-element group 610:  transition  input  no-bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	604 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	66 
    -- CP-element group 610:  members (4) 
      -- CP-element group 610: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/$exit
      -- CP-element group 610: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_update_completed_
      -- CP-element group 610: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Update/$exit
      -- CP-element group 610: 	 branch_block_stmt_1353/assign_stmt_2206_to_assign_stmt_2216/SLT_f64_u1_2215_Update/ca
      -- 
    ca_10264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 610_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_f64_u1_2215_inst_ack_1, ack => minSumDecode_CP_6680_elements(610)); -- 
    -- CP-element group 611:  transition  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	66 
    -- CP-element group 611: successors 
    -- CP-element group 611:  members (1) 
      -- CP-element group 611: 	 branch_block_stmt_1353/if_stmt_2217_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(611) <= minSumDecode_CP_6680_elements(66);
    -- CP-element group 612:  transition  output  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	66 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	613 
    -- CP-element group 612:  members (3) 
      -- CP-element group 612: 	 branch_block_stmt_1353/if_stmt_2217_eval_test/$entry
      -- CP-element group 612: 	 branch_block_stmt_1353/if_stmt_2217_eval_test/$exit
      -- CP-element group 612: 	 branch_block_stmt_1353/if_stmt_2217_eval_test/branch_req
      -- 
    branch_req_10272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(612), ack => if_stmt_2217_branch_req_0); -- 
    minSumDecode_CP_6680_elements(612) <= minSumDecode_CP_6680_elements(66);
    -- CP-element group 613:  branch  place  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	612 
    -- CP-element group 613: successors 
    -- CP-element group 613: 	614 
    -- CP-element group 613: 	616 
    -- CP-element group 613:  members (1) 
      -- CP-element group 613: 	 branch_block_stmt_1353/R_iNsTr_123_2218_place
      -- 
    minSumDecode_CP_6680_elements(613) <= minSumDecode_CP_6680_elements(612);
    -- CP-element group 614:  transition  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	613 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	615 
    -- CP-element group 614:  members (1) 
      -- CP-element group 614: 	 branch_block_stmt_1353/if_stmt_2217_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(614) <= minSumDecode_CP_6680_elements(613);
    -- CP-element group 615:  transition  input  no-bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	614 
    -- CP-element group 615: successors 
    -- CP-element group 615: 	618 
    -- CP-element group 615:  members (2) 
      -- CP-element group 615: 	 branch_block_stmt_1353/if_stmt_2217_if_link/$exit
      -- CP-element group 615: 	 branch_block_stmt_1353/if_stmt_2217_if_link/if_choice_transition
      -- 
    if_choice_transition_10277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2217_branch_ack_1, ack => minSumDecode_CP_6680_elements(615)); -- 
    -- CP-element group 616:  transition  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	613 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	617 
    -- CP-element group 616:  members (1) 
      -- CP-element group 616: 	 branch_block_stmt_1353/if_stmt_2217_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(616) <= minSumDecode_CP_6680_elements(613);
    -- CP-element group 617:  transition  input  no-bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	616 
    -- CP-element group 617: successors 
    -- CP-element group 617: 	619 
    -- CP-element group 617:  members (2) 
      -- CP-element group 617: 	 branch_block_stmt_1353/if_stmt_2217_else_link/$exit
      -- CP-element group 617: 	 branch_block_stmt_1353/if_stmt_2217_else_link/else_choice_transition
      -- 
    else_choice_transition_10281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2217_branch_ack_0, ack => minSumDecode_CP_6680_elements(617)); -- 
    -- CP-element group 618:  place  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	615 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	1073 
    -- CP-element group 618:  members (1) 
      -- CP-element group 618: 	 branch_block_stmt_1353/bb_34_bb_35
      -- 
    minSumDecode_CP_6680_elements(618) <= minSumDecode_CP_6680_elements(615);
    -- CP-element group 619:  place  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	617 
    -- CP-element group 619: successors 
    -- CP-element group 619: 	1076 
    -- CP-element group 619:  members (1) 
      -- CP-element group 619: 	 branch_block_stmt_1353/bb_34_bb_36
      -- 
    minSumDecode_CP_6680_elements(619) <= minSumDecode_CP_6680_elements(617);
    -- CP-element group 620:  fork  transition  output  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	67 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	621 
    -- CP-element group 620: 	622 
    -- CP-element group 620:  members (17) 
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_update_start_
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/STORE_is_decoded_2224_Split/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/STORE_is_decoded_2224_Split/$exit
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/STORE_is_decoded_2224_Split/split_req
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/STORE_is_decoded_2224_Split/split_ack
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/word_0/cr
      -- 
    cr_10318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(620), ack => STORE_is_decoded_2224_store_0_req_1); -- 
    rr_10307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(620), ack => STORE_is_decoded_2224_store_0_req_0); -- 
    minSumDecode_CP_6680_elements(620) <= minSumDecode_CP_6680_elements(67);
    -- CP-element group 621:  transition  input  no-bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	620 
    -- CP-element group 621: successors 
    -- CP-element group 621:  members (5) 
      -- CP-element group 621: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_sample_completed_
      -- CP-element group 621: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/$exit
      -- CP-element group 621: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/$exit
      -- CP-element group 621: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/word_0/$exit
      -- CP-element group 621: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Sample/word_access_start/word_0/ra
      -- 
    ra_10308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2224_store_0_ack_0, ack => minSumDecode_CP_6680_elements(621)); -- 
    -- CP-element group 622:  transition  input  no-bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	620 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	68 
    -- CP-element group 622:  members (6) 
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/$exit
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_update_completed_
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/$exit
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/$exit
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/word_0/$exit
      -- CP-element group 622: 	 branch_block_stmt_1353/assign_stmt_2227/STORE_is_decoded_2224_Update/word_access_complete/word_0/ca
      -- 
    ca_10319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_is_decoded_2224_store_0_ack_1, ack => minSumDecode_CP_6680_elements(622)); -- 
    -- CP-element group 623:  join  fork  transition  output  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	69 
    -- CP-element group 623: successors 
    -- CP-element group 623: 	624 
    -- CP-element group 623: 	625 
    -- CP-element group 623:  members (31) 
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_sample_start_
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_update_start_
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_address_calculated
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_word_address_calculated
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_root_address_calculated
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_address_resized
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_addr_resize/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_addr_resize/$exit
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_addr_resize/base_resize_req
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_addr_resize/base_resize_ack
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_plus_offset/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_plus_offset/$exit
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_plus_offset/sum_rename_req
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_base_plus_offset/sum_rename_ack
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_word_addrgen/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_word_addrgen/$exit
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_word_addrgen/root_register_req
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_word_addrgen/root_register_ack
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/ptr_deref_2239_Split/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/ptr_deref_2239_Split/$exit
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/ptr_deref_2239_Split/split_req
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/ptr_deref_2239_Split/split_ack
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/word_0/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/word_0/rr
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/word_0/$entry
      -- CP-element group 623: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/word_0/cr
      -- 
    cr_10371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(623), ack => ptr_deref_2239_store_0_req_1); -- 
    rr_10360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(623), ack => ptr_deref_2239_store_0_req_0); -- 
    minSumDecode_CP_6680_elements(623) <= minSumDecode_CP_6680_elements(69);
    -- CP-element group 624:  transition  input  no-bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	623 
    -- CP-element group 624: successors 
    -- CP-element group 624:  members (5) 
      -- CP-element group 624: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_sample_completed_
      -- CP-element group 624: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/$exit
      -- CP-element group 624: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/$exit
      -- CP-element group 624: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/word_0/$exit
      -- CP-element group 624: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Sample/word_access_start/word_0/ra
      -- 
    ra_10361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2239_store_0_ack_0, ack => minSumDecode_CP_6680_elements(624)); -- 
    -- CP-element group 625:  transition  input  no-bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	623 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	70 
    -- CP-element group 625:  members (6) 
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/$exit
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_update_completed_
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/$exit
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/$exit
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/word_0/$exit
      -- CP-element group 625: 	 branch_block_stmt_1353/assign_stmt_2242/ptr_deref_2239_Update/word_access_complete/word_0/ca
      -- 
    ca_10372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2239_store_0_ack_1, ack => minSumDecode_CP_6680_elements(625)); -- 
    -- CP-element group 626:  fork  transition  output  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	71 
    -- CP-element group 626: successors 
    -- CP-element group 626: 	627 
    -- CP-element group 626: 	628 
    -- CP-element group 626: 	630 
    -- CP-element group 626:  members (10) 
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/$entry
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_sample_start_
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_update_start_
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Sample/$entry
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Sample/rr
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Update/$entry
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Update/cr
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_update_start_
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Update/$entry
      -- CP-element group 626: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Update/cr
      -- 
    rr_10383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(626), ack => ADD_u64_u64_2258_inst_req_0); -- 
    cr_10388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(626), ack => ADD_u64_u64_2258_inst_req_1); -- 
    cr_10402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(626), ack => EQ_u64_u1_2263_inst_req_1); -- 
    minSumDecode_CP_6680_elements(626) <= minSumDecode_CP_6680_elements(71);
    -- CP-element group 627:  transition  input  no-bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	626 
    -- CP-element group 627: successors 
    -- CP-element group 627:  members (3) 
      -- CP-element group 627: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_sample_completed_
      -- CP-element group 627: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Sample/$exit
      -- CP-element group 627: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Sample/ra
      -- 
    ra_10384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2258_inst_ack_0, ack => minSumDecode_CP_6680_elements(627)); -- 
    -- CP-element group 628:  transition  input  output  no-bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	626 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	629 
    -- CP-element group 628:  members (6) 
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_update_completed_
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Update/$exit
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/ADD_u64_u64_2258_Update/ca
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_sample_start_
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Sample/$entry
      -- CP-element group 628: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Sample/rr
      -- 
    ca_10389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2258_inst_ack_1, ack => minSumDecode_CP_6680_elements(628)); -- 
    rr_10397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(628), ack => EQ_u64_u1_2263_inst_req_0); -- 
    -- CP-element group 629:  transition  input  no-bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	628 
    -- CP-element group 629: successors 
    -- CP-element group 629:  members (3) 
      -- CP-element group 629: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_sample_completed_
      -- CP-element group 629: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Sample/$exit
      -- CP-element group 629: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Sample/ra
      -- 
    ra_10398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2263_inst_ack_0, ack => minSumDecode_CP_6680_elements(629)); -- 
    -- CP-element group 630:  transition  input  no-bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	626 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	72 
    -- CP-element group 630:  members (4) 
      -- CP-element group 630: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/$exit
      -- CP-element group 630: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_update_completed_
      -- CP-element group 630: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Update/$exit
      -- CP-element group 630: 	 branch_block_stmt_1353/assign_stmt_2259_to_assign_stmt_2264/EQ_u64_u1_2263_Update/ca
      -- 
    ca_10403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2263_inst_ack_1, ack => minSumDecode_CP_6680_elements(630)); -- 
    -- CP-element group 631:  transition  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	72 
    -- CP-element group 631: successors 
    -- CP-element group 631:  members (1) 
      -- CP-element group 631: 	 branch_block_stmt_1353/if_stmt_2265_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(631) <= minSumDecode_CP_6680_elements(72);
    -- CP-element group 632:  transition  output  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	72 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	633 
    -- CP-element group 632:  members (3) 
      -- CP-element group 632: 	 branch_block_stmt_1353/if_stmt_2265_eval_test/$entry
      -- CP-element group 632: 	 branch_block_stmt_1353/if_stmt_2265_eval_test/$exit
      -- CP-element group 632: 	 branch_block_stmt_1353/if_stmt_2265_eval_test/branch_req
      -- 
    branch_req_10411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(632), ack => if_stmt_2265_branch_req_0); -- 
    minSumDecode_CP_6680_elements(632) <= minSumDecode_CP_6680_elements(72);
    -- CP-element group 633:  branch  place  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	632 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	634 
    -- CP-element group 633: 	636 
    -- CP-element group 633:  members (1) 
      -- CP-element group 633: 	 branch_block_stmt_1353/R_exitcond16_2266_place
      -- 
    minSumDecode_CP_6680_elements(633) <= minSumDecode_CP_6680_elements(632);
    -- CP-element group 634:  transition  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	633 
    -- CP-element group 634: successors 
    -- CP-element group 634: 	635 
    -- CP-element group 634:  members (1) 
      -- CP-element group 634: 	 branch_block_stmt_1353/if_stmt_2265_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(634) <= minSumDecode_CP_6680_elements(633);
    -- CP-element group 635:  transition  input  no-bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	634 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	638 
    -- CP-element group 635:  members (2) 
      -- CP-element group 635: 	 branch_block_stmt_1353/if_stmt_2265_if_link/$exit
      -- CP-element group 635: 	 branch_block_stmt_1353/if_stmt_2265_if_link/if_choice_transition
      -- 
    if_choice_transition_10416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2265_branch_ack_1, ack => minSumDecode_CP_6680_elements(635)); -- 
    -- CP-element group 636:  transition  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	633 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	637 
    -- CP-element group 636:  members (1) 
      -- CP-element group 636: 	 branch_block_stmt_1353/if_stmt_2265_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(636) <= minSumDecode_CP_6680_elements(633);
    -- CP-element group 637:  transition  input  no-bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	636 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	639 
    -- CP-element group 637:  members (2) 
      -- CP-element group 637: 	 branch_block_stmt_1353/if_stmt_2265_else_link/$exit
      -- CP-element group 637: 	 branch_block_stmt_1353/if_stmt_2265_else_link/else_choice_transition
      -- 
    else_choice_transition_10420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2265_branch_ack_0, ack => minSumDecode_CP_6680_elements(637)); -- 
    -- CP-element group 638:  place  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	635 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	1101 
    -- CP-element group 638:  members (1) 
      -- CP-element group 638: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit
      -- 
    minSumDecode_CP_6680_elements(638) <= minSumDecode_CP_6680_elements(635);
    -- CP-element group 639:  place  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	637 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	1032 
    -- CP-element group 639:  members (1) 
      -- CP-element group 639: 	 branch_block_stmt_1353/bb_37_bb_29
      -- 
    minSumDecode_CP_6680_elements(639) <= minSumDecode_CP_6680_elements(637);
    -- CP-element group 640:  fork  transition  output  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	73 
    -- CP-element group 640: successors 
    -- CP-element group 640: 	641 
    -- CP-element group 640: 	642 
    -- CP-element group 640:  members (7) 
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/$entry
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_sample_start_
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_update_start_
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Sample/$entry
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Sample/rr
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Update/$entry
      -- CP-element group 640: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Update/cr
      -- 
    rr_10433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(640), ack => EQ_u16_u1_2281_inst_req_0); -- 
    cr_10438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(640), ack => EQ_u16_u1_2281_inst_req_1); -- 
    minSumDecode_CP_6680_elements(640) <= minSumDecode_CP_6680_elements(73);
    -- CP-element group 641:  transition  input  no-bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	640 
    -- CP-element group 641: successors 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_sample_completed_
      -- CP-element group 641: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Sample/$exit
      -- CP-element group 641: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Sample/ra
      -- 
    ra_10434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 641_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2281_inst_ack_0, ack => minSumDecode_CP_6680_elements(641)); -- 
    -- CP-element group 642:  transition  input  no-bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	640 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	74 
    -- CP-element group 642:  members (4) 
      -- CP-element group 642: 	 branch_block_stmt_1353/assign_stmt_2282/$exit
      -- CP-element group 642: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_update_completed_
      -- CP-element group 642: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Update/$exit
      -- CP-element group 642: 	 branch_block_stmt_1353/assign_stmt_2282/EQ_u16_u1_2281_Update/ca
      -- 
    ca_10439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 642_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2281_inst_ack_1, ack => minSumDecode_CP_6680_elements(642)); -- 
    -- CP-element group 643:  transition  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	74 
    -- CP-element group 643: successors 
    -- CP-element group 643:  members (1) 
      -- CP-element group 643: 	 branch_block_stmt_1353/if_stmt_2283_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(643) <= minSumDecode_CP_6680_elements(74);
    -- CP-element group 644:  transition  output  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	74 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644:  members (3) 
      -- CP-element group 644: 	 branch_block_stmt_1353/if_stmt_2283_eval_test/$entry
      -- CP-element group 644: 	 branch_block_stmt_1353/if_stmt_2283_eval_test/$exit
      -- CP-element group 644: 	 branch_block_stmt_1353/if_stmt_2283_eval_test/branch_req
      -- 
    branch_req_10447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(644), ack => if_stmt_2283_branch_req_0); -- 
    minSumDecode_CP_6680_elements(644) <= minSumDecode_CP_6680_elements(74);
    -- CP-element group 645:  branch  place  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	646 
    -- CP-element group 645: 	648 
    -- CP-element group 645:  members (1) 
      -- CP-element group 645: 	 branch_block_stmt_1353/R_iNsTr_130_2284_place
      -- 
    minSumDecode_CP_6680_elements(645) <= minSumDecode_CP_6680_elements(644);
    -- CP-element group 646:  transition  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	645 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646:  members (1) 
      -- CP-element group 646: 	 branch_block_stmt_1353/if_stmt_2283_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(646) <= minSumDecode_CP_6680_elements(645);
    -- CP-element group 647:  transition  input  no-bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	650 
    -- CP-element group 647:  members (2) 
      -- CP-element group 647: 	 branch_block_stmt_1353/if_stmt_2283_if_link/$exit
      -- CP-element group 647: 	 branch_block_stmt_1353/if_stmt_2283_if_link/if_choice_transition
      -- 
    if_choice_transition_10452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2283_branch_ack_1, ack => minSumDecode_CP_6680_elements(647)); -- 
    -- CP-element group 648:  transition  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	645 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (1) 
      -- CP-element group 648: 	 branch_block_stmt_1353/if_stmt_2283_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(648) <= minSumDecode_CP_6680_elements(645);
    -- CP-element group 649:  transition  input  no-bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649: 	651 
    -- CP-element group 649:  members (2) 
      -- CP-element group 649: 	 branch_block_stmt_1353/if_stmt_2283_else_link/$exit
      -- CP-element group 649: 	 branch_block_stmt_1353/if_stmt_2283_else_link/else_choice_transition
      -- 
    else_choice_transition_10456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2283_branch_ack_0, ack => minSumDecode_CP_6680_elements(649)); -- 
    -- CP-element group 650:  place  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	647 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	1178 
    -- CP-element group 650:  members (1) 
      -- CP-element group 650: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread
      -- 
    minSumDecode_CP_6680_elements(650) <= minSumDecode_CP_6680_elements(647);
    -- CP-element group 651:  place  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	649 
    -- CP-element group 651: successors 
    -- CP-element group 651: 	1108 
    -- CP-element group 651:  members (1) 
      -- CP-element group 651: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_bb_39
      -- 
    minSumDecode_CP_6680_elements(651) <= minSumDecode_CP_6680_elements(649);
    -- CP-element group 652:  fork  transition  output  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	75 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	653 
    -- CP-element group 652: 	654 
    -- CP-element group 652: 	656 
    -- CP-element group 652:  members (16) 
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_sample_start_
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_update_start_
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_word_address_calculated
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_root_address_calculated
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/word_0/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/word_0/rr
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/word_0/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/word_0/cr
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_update_start_
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Update/$entry
      -- CP-element group 652: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Update/cr
      -- 
    cr_10488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(652), ack => LOAD_nrows_2291_load_0_req_1); -- 
    rr_10477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(652), ack => LOAD_nrows_2291_load_0_req_0); -- 
    cr_10507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(652), ack => EQ_u16_u1_2297_inst_req_1); -- 
    minSumDecode_CP_6680_elements(652) <= minSumDecode_CP_6680_elements(75);
    -- CP-element group 653:  transition  input  no-bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	652 
    -- CP-element group 653: successors 
    -- CP-element group 653:  members (5) 
      -- CP-element group 653: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_sample_completed_
      -- CP-element group 653: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/$exit
      -- CP-element group 653: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/$exit
      -- CP-element group 653: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/word_0/$exit
      -- CP-element group 653: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Sample/word_access_start/word_0/ra
      -- 
    ra_10478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 653_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_2291_load_0_ack_0, ack => minSumDecode_CP_6680_elements(653)); -- 
    -- CP-element group 654:  transition  input  output  no-bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	652 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	655 
    -- CP-element group 654:  members (12) 
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_update_completed_
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/$exit
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/$exit
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/word_0/$exit
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/word_access_complete/word_0/ca
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/LOAD_nrows_2291_Merge/$entry
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/LOAD_nrows_2291_Merge/$exit
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/LOAD_nrows_2291_Merge/merge_req
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/LOAD_nrows_2291_Update/LOAD_nrows_2291_Merge/merge_ack
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_sample_start_
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Sample/$entry
      -- CP-element group 654: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Sample/rr
      -- 
    ca_10489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 654_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_nrows_2291_load_0_ack_1, ack => minSumDecode_CP_6680_elements(654)); -- 
    rr_10502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(654), ack => EQ_u16_u1_2297_inst_req_0); -- 
    -- CP-element group 655:  transition  input  no-bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	654 
    -- CP-element group 655: successors 
    -- CP-element group 655:  members (3) 
      -- CP-element group 655: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_sample_completed_
      -- CP-element group 655: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Sample/$exit
      -- CP-element group 655: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Sample/ra
      -- 
    ra_10503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2297_inst_ack_0, ack => minSumDecode_CP_6680_elements(655)); -- 
    -- CP-element group 656:  transition  input  no-bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	652 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	76 
    -- CP-element group 656:  members (4) 
      -- CP-element group 656: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/$exit
      -- CP-element group 656: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_update_completed_
      -- CP-element group 656: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Update/$exit
      -- CP-element group 656: 	 branch_block_stmt_1353/assign_stmt_2292_to_assign_stmt_2298/EQ_u16_u1_2297_Update/ca
      -- 
    ca_10508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2297_inst_ack_1, ack => minSumDecode_CP_6680_elements(656)); -- 
    -- CP-element group 657:  transition  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	76 
    -- CP-element group 657: successors 
    -- CP-element group 657:  members (1) 
      -- CP-element group 657: 	 branch_block_stmt_1353/if_stmt_2299_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(657) <= minSumDecode_CP_6680_elements(76);
    -- CP-element group 658:  transition  output  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	76 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (3) 
      -- CP-element group 658: 	 branch_block_stmt_1353/if_stmt_2299_eval_test/$entry
      -- CP-element group 658: 	 branch_block_stmt_1353/if_stmt_2299_eval_test/$exit
      -- CP-element group 658: 	 branch_block_stmt_1353/if_stmt_2299_eval_test/branch_req
      -- 
    branch_req_10516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(658), ack => if_stmt_2299_branch_req_0); -- 
    minSumDecode_CP_6680_elements(658) <= minSumDecode_CP_6680_elements(76);
    -- CP-element group 659:  branch  place  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	660 
    -- CP-element group 659: 	662 
    -- CP-element group 659:  members (1) 
      -- CP-element group 659: 	 branch_block_stmt_1353/R_iNsTr_133_2300_place
      -- 
    minSumDecode_CP_6680_elements(659) <= minSumDecode_CP_6680_elements(658);
    -- CP-element group 660:  transition  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	659 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	661 
    -- CP-element group 660:  members (1) 
      -- CP-element group 660: 	 branch_block_stmt_1353/if_stmt_2299_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(660) <= minSumDecode_CP_6680_elements(659);
    -- CP-element group 661:  transition  input  no-bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	660 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	664 
    -- CP-element group 661:  members (2) 
      -- CP-element group 661: 	 branch_block_stmt_1353/if_stmt_2299_if_link/$exit
      -- CP-element group 661: 	 branch_block_stmt_1353/if_stmt_2299_if_link/if_choice_transition
      -- 
    if_choice_transition_10521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2299_branch_ack_1, ack => minSumDecode_CP_6680_elements(661)); -- 
    -- CP-element group 662:  transition  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	659 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	663 
    -- CP-element group 662:  members (1) 
      -- CP-element group 662: 	 branch_block_stmt_1353/if_stmt_2299_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(662) <= minSumDecode_CP_6680_elements(659);
    -- CP-element group 663:  transition  input  no-bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	662 
    -- CP-element group 663: successors 
    -- CP-element group 663: 	665 
    -- CP-element group 663:  members (2) 
      -- CP-element group 663: 	 branch_block_stmt_1353/if_stmt_2299_else_link/$exit
      -- CP-element group 663: 	 branch_block_stmt_1353/if_stmt_2299_else_link/else_choice_transition
      -- 
    else_choice_transition_10525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2299_branch_ack_0, ack => minSumDecode_CP_6680_elements(663)); -- 
    -- CP-element group 664:  place  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	661 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	1174 
    -- CP-element group 664:  members (1) 
      -- CP-element group 664: 	 branch_block_stmt_1353/bb_39_updateMessagex_xexit
      -- 
    minSumDecode_CP_6680_elements(664) <= minSumDecode_CP_6680_elements(661);
    -- CP-element group 665:  place  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	663 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	1111 
    -- CP-element group 665:  members (1) 
      -- CP-element group 665: 	 branch_block_stmt_1353/bb_39_bbx_xnph4x_xi
      -- 
    minSumDecode_CP_6680_elements(665) <= minSumDecode_CP_6680_elements(663);
    -- CP-element group 666:  fork  transition  output  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	77 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	667 
    -- CP-element group 666: 	668 
    -- CP-element group 666: 	670 
    -- CP-element group 666: 	671 
    -- CP-element group 666: 	672 
    -- CP-element group 666: 	673 
    -- CP-element group 666: 	674 
    -- CP-element group 666: 	676 
    -- CP-element group 666: 	678 
    -- CP-element group 666: 	681 
    -- CP-element group 666: 	682 
    -- CP-element group 666: 	683 
    -- CP-element group 666: 	684 
    -- CP-element group 666: 	685 
    -- CP-element group 666: 	687 
    -- CP-element group 666: 	689 
    -- CP-element group 666:  members (49) 
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_complete/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_complete/req
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_update_start_
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_update_start_
      -- 
    rr_10538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => type_cast_2308_inst_req_0); -- 
    cr_10543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => type_cast_2308_inst_req_1); -- 
    cr_10557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u32_u32_2314_inst_req_1); -- 
    rr_10566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => UGT_u16_u1_2320_inst_req_0); -- 
    cr_10571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => UGT_u16_u1_2320_inst_req_1); -- 
    rr_10580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u16_u16_2326_inst_req_0); -- 
    cr_10585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u16_u16_2326_inst_req_1); -- 
    cr_10599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => type_cast_2330_inst_req_1); -- 
    cr_10613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u64_u64_2336_inst_req_1); -- 
    req_10627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => MUX_2343_inst_req_1); -- 
    rr_10636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u16_u16_2349_inst_req_0); -- 
    cr_10641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u16_u16_2349_inst_req_1); -- 
    rr_10650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => type_cast_2353_inst_req_0); -- 
    cr_10655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => type_cast_2353_inst_req_1); -- 
    cr_10669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u64_u64_2359_inst_req_1); -- 
    cr_10683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(666), ack => ADD_u64_u64_2365_inst_req_1); -- 
    minSumDecode_CP_6680_elements(666) <= minSumDecode_CP_6680_elements(77);
    -- CP-element group 667:  transition  input  no-bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	666 
    -- CP-element group 667: successors 
    -- CP-element group 667:  members (3) 
      -- CP-element group 667: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_sample_completed_
      -- CP-element group 667: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Sample/$exit
      -- CP-element group 667: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Sample/ra
      -- 
    ra_10539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_0, ack => minSumDecode_CP_6680_elements(667)); -- 
    -- CP-element group 668:  transition  input  output  no-bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	666 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	669 
    -- CP-element group 668:  members (6) 
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_update_completed_
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Update/$exit
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2308_Update/ca
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_sample_start_
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Sample/$entry
      -- CP-element group 668: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Sample/rr
      -- 
    ca_10544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 668_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_1, ack => minSumDecode_CP_6680_elements(668)); -- 
    rr_10552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(668), ack => ADD_u32_u32_2314_inst_req_0); -- 
    -- CP-element group 669:  transition  input  no-bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	668 
    -- CP-element group 669: successors 
    -- CP-element group 669:  members (3) 
      -- CP-element group 669: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_sample_completed_
      -- CP-element group 669: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Sample/$exit
      -- CP-element group 669: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Sample/ra
      -- 
    ra_10553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2314_inst_ack_0, ack => minSumDecode_CP_6680_elements(669)); -- 
    -- CP-element group 670:  transition  input  no-bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	666 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	690 
    -- CP-element group 670:  members (3) 
      -- CP-element group 670: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_update_completed_
      -- CP-element group 670: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Update/$exit
      -- CP-element group 670: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u32_u32_2314_Update/ca
      -- 
    ca_10558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 670_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2314_inst_ack_1, ack => minSumDecode_CP_6680_elements(670)); -- 
    -- CP-element group 671:  transition  input  no-bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	666 
    -- CP-element group 671: successors 
    -- CP-element group 671:  members (3) 
      -- CP-element group 671: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_sample_completed_
      -- CP-element group 671: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Sample/$exit
      -- CP-element group 671: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Sample/ra
      -- 
    ra_10567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_2320_inst_ack_0, ack => minSumDecode_CP_6680_elements(671)); -- 
    -- CP-element group 672:  transition  input  no-bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	666 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	679 
    -- CP-element group 672:  members (3) 
      -- CP-element group 672: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_update_completed_
      -- CP-element group 672: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Update/$exit
      -- CP-element group 672: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/UGT_u16_u1_2320_Update/ca
      -- 
    ca_10572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UGT_u16_u1_2320_inst_ack_1, ack => minSumDecode_CP_6680_elements(672)); -- 
    -- CP-element group 673:  transition  input  no-bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	666 
    -- CP-element group 673: successors 
    -- CP-element group 673:  members (3) 
      -- CP-element group 673: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_sample_completed_
      -- CP-element group 673: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Sample/$exit
      -- CP-element group 673: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Sample/ra
      -- 
    ra_10581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 673_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2326_inst_ack_0, ack => minSumDecode_CP_6680_elements(673)); -- 
    -- CP-element group 674:  transition  input  output  no-bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	666 
    -- CP-element group 674: successors 
    -- CP-element group 674: 	675 
    -- CP-element group 674:  members (6) 
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_update_completed_
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Update/$exit
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2326_Update/ca
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Sample/rr
      -- 
    ca_10586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 674_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2326_inst_ack_1, ack => minSumDecode_CP_6680_elements(674)); -- 
    rr_10594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(674), ack => type_cast_2330_inst_req_0); -- 
    -- CP-element group 675:  transition  input  no-bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	674 
    -- CP-element group 675: successors 
    -- CP-element group 675:  members (3) 
      -- CP-element group 675: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_sample_completed_
      -- CP-element group 675: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Sample/$exit
      -- CP-element group 675: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Sample/ra
      -- 
    ra_10595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2330_inst_ack_0, ack => minSumDecode_CP_6680_elements(675)); -- 
    -- CP-element group 676:  transition  input  output  no-bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	666 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	677 
    -- CP-element group 676:  members (6) 
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_update_completed_
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Update/$exit
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2330_Update/ca
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_sample_start_
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Sample/$entry
      -- CP-element group 676: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Sample/rr
      -- 
    ca_10600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2330_inst_ack_1, ack => minSumDecode_CP_6680_elements(676)); -- 
    rr_10608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(676), ack => ADD_u64_u64_2336_inst_req_0); -- 
    -- CP-element group 677:  transition  input  no-bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	676 
    -- CP-element group 677: successors 
    -- CP-element group 677:  members (3) 
      -- CP-element group 677: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_sample_completed_
      -- CP-element group 677: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Sample/$exit
      -- CP-element group 677: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Sample/ra
      -- 
    ra_10609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 677_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2336_inst_ack_0, ack => minSumDecode_CP_6680_elements(677)); -- 
    -- CP-element group 678:  transition  input  no-bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	666 
    -- CP-element group 678: successors 
    -- CP-element group 678: 	679 
    -- CP-element group 678:  members (3) 
      -- CP-element group 678: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_update_completed_
      -- CP-element group 678: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Update/$exit
      -- CP-element group 678: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2336_Update/ca
      -- 
    ca_10614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2336_inst_ack_1, ack => minSumDecode_CP_6680_elements(678)); -- 
    -- CP-element group 679:  join  transition  output  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	672 
    -- CP-element group 679: 	678 
    -- CP-element group 679: successors 
    -- CP-element group 679: 	680 
    -- CP-element group 679:  members (3) 
      -- CP-element group 679: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_sample_start_
      -- CP-element group 679: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_start/$entry
      -- CP-element group 679: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_start/req
      -- 
    req_10622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(679), ack => MUX_2343_inst_req_0); -- 
    minSumDecode_cp_element_group_679: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_679"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(672) & minSumDecode_CP_6680_elements(678);
      gj_minSumDecode_cp_element_group_679 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(679), clk => clk, reset => reset); --
    end block;
    -- CP-element group 680:  transition  input  no-bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	679 
    -- CP-element group 680: successors 
    -- CP-element group 680: 	690 
    -- CP-element group 680:  members (3) 
      -- CP-element group 680: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_sample_completed_
      -- CP-element group 680: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_start/$exit
      -- CP-element group 680: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_start/ack
      -- 
    ack_10623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2343_inst_ack_0, ack => minSumDecode_CP_6680_elements(680)); -- 
    -- CP-element group 681:  transition  input  no-bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	666 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	690 
    -- CP-element group 681:  members (3) 
      -- CP-element group 681: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_update_completed_
      -- CP-element group 681: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_complete/$exit
      -- CP-element group 681: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/MUX_2343_complete/ack
      -- 
    ack_10628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2343_inst_ack_1, ack => minSumDecode_CP_6680_elements(681)); -- 
    -- CP-element group 682:  transition  input  no-bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	666 
    -- CP-element group 682: successors 
    -- CP-element group 682:  members (3) 
      -- CP-element group 682: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_sample_completed_
      -- CP-element group 682: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Sample/$exit
      -- CP-element group 682: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Sample/ra
      -- 
    ra_10637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 682_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2349_inst_ack_0, ack => minSumDecode_CP_6680_elements(682)); -- 
    -- CP-element group 683:  transition  input  no-bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	666 
    -- CP-element group 683: successors 
    -- CP-element group 683: 	690 
    -- CP-element group 683:  members (3) 
      -- CP-element group 683: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_update_completed_
      -- CP-element group 683: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Update/$exit
      -- CP-element group 683: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u16_u16_2349_Update/ca
      -- 
    ca_10642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2349_inst_ack_1, ack => minSumDecode_CP_6680_elements(683)); -- 
    -- CP-element group 684:  transition  input  no-bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	666 
    -- CP-element group 684: successors 
    -- CP-element group 684:  members (3) 
      -- CP-element group 684: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_sample_completed_
      -- CP-element group 684: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Sample/$exit
      -- CP-element group 684: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Sample/ra
      -- 
    ra_10651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 684_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_0, ack => minSumDecode_CP_6680_elements(684)); -- 
    -- CP-element group 685:  fork  transition  input  output  no-bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	666 
    -- CP-element group 685: successors 
    -- CP-element group 685: 	686 
    -- CP-element group 685: 	688 
    -- CP-element group 685:  members (9) 
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_update_completed_
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Update/$exit
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/type_cast_2353_Update/ca
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_sample_start_
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Sample/$entry
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Sample/rr
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_sample_start_
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Sample/$entry
      -- CP-element group 685: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Sample/rr
      -- 
    ca_10656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 685_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_1, ack => minSumDecode_CP_6680_elements(685)); -- 
    rr_10664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(685), ack => ADD_u64_u64_2359_inst_req_0); -- 
    rr_10678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(685), ack => ADD_u64_u64_2365_inst_req_0); -- 
    -- CP-element group 686:  transition  input  no-bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	685 
    -- CP-element group 686: successors 
    -- CP-element group 686:  members (3) 
      -- CP-element group 686: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_sample_completed_
      -- CP-element group 686: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Sample/$exit
      -- CP-element group 686: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Sample/ra
      -- 
    ra_10665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2359_inst_ack_0, ack => minSumDecode_CP_6680_elements(686)); -- 
    -- CP-element group 687:  transition  input  no-bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	666 
    -- CP-element group 687: successors 
    -- CP-element group 687: 	690 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_update_completed_
      -- CP-element group 687: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Update/$exit
      -- CP-element group 687: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2359_Update/ca
      -- 
    ca_10670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2359_inst_ack_1, ack => minSumDecode_CP_6680_elements(687)); -- 
    -- CP-element group 688:  transition  input  no-bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	685 
    -- CP-element group 688: successors 
    -- CP-element group 688:  members (3) 
      -- CP-element group 688: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_sample_completed_
      -- CP-element group 688: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Sample/$exit
      -- CP-element group 688: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Sample/ra
      -- 
    ra_10679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2365_inst_ack_0, ack => minSumDecode_CP_6680_elements(688)); -- 
    -- CP-element group 689:  transition  input  no-bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	666 
    -- CP-element group 689: successors 
    -- CP-element group 689: 	690 
    -- CP-element group 689:  members (3) 
      -- CP-element group 689: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Update/ca
      -- CP-element group 689: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_Update/$exit
      -- CP-element group 689: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/ADD_u64_u64_2365_update_completed_
      -- 
    ca_10684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 689_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2365_inst_ack_1, ack => minSumDecode_CP_6680_elements(689)); -- 
    -- CP-element group 690:  join  transition  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	670 
    -- CP-element group 690: 	680 
    -- CP-element group 690: 	681 
    -- CP-element group 690: 	683 
    -- CP-element group 690: 	687 
    -- CP-element group 690: 	689 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	78 
    -- CP-element group 690:  members (1) 
      -- CP-element group 690: 	 branch_block_stmt_1353/assign_stmt_2309_to_assign_stmt_2366/$exit
      -- 
    minSumDecode_cp_element_group_690: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_690"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(670) & minSumDecode_CP_6680_elements(680) & minSumDecode_CP_6680_elements(681) & minSumDecode_CP_6680_elements(683) & minSumDecode_CP_6680_elements(687) & minSumDecode_CP_6680_elements(689);
      gj_minSumDecode_cp_element_group_690 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(690), clk => clk, reset => reset); --
    end block;
    -- CP-element group 691:  fork  transition  output  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	79 
    -- CP-element group 691: successors 
    -- CP-element group 691: 	692 
    -- CP-element group 691: 	693 
    -- CP-element group 691: 	695 
    -- CP-element group 691: 	696 
    -- CP-element group 691: 	697 
    -- CP-element group 691: 	698 
    -- CP-element group 691: 	699 
    -- CP-element group 691: 	701 
    -- CP-element group 691: 	703 
    -- CP-element group 691:  members (28) 
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Sample/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Sample/rr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Update/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Sample/rr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Update/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Update/cr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Update/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Update/cr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_sample_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Sample/rr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_complete/req
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Sample/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_complete/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_sample_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Sample/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_sample_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Update/cr
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_complete/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_complete/req
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_update_start_
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Update/$entry
      -- CP-element group 691: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Update/cr
      -- 
    rr_10695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => ADD_u64_u64_2380_inst_req_0); -- 
    cr_10700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => ADD_u64_u64_2380_inst_req_1); -- 
    req_10739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => addr_of_2385_final_reg_req_1); -- 
    rr_10748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => type_cast_2389_inst_req_0); -- 
    cr_10753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => type_cast_2389_inst_req_1); -- 
    rr_10762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => ADD_u64_u64_2394_inst_req_0); -- 
    cr_10767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => ADD_u64_u64_2394_inst_req_1); -- 
    req_10806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => addr_of_2399_final_reg_req_1); -- 
    cr_10820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(691), ack => EQ_u32_u1_2404_inst_req_1); -- 
    minSumDecode_CP_6680_elements(691) <= minSumDecode_CP_6680_elements(79);
    -- CP-element group 692:  transition  input  no-bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	691 
    -- CP-element group 692: successors 
    -- CP-element group 692:  members (3) 
      -- CP-element group 692: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Sample/ra
      -- CP-element group 692: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Sample/$exit
      -- CP-element group 692: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_sample_completed_
      -- 
    ra_10696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2380_inst_ack_0, ack => minSumDecode_CP_6680_elements(692)); -- 
    -- CP-element group 693:  transition  input  output  no-bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	691 
    -- CP-element group 693: successors 
    -- CP-element group 693: 	694 
    -- CP-element group 693:  members (27) 
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Update/ca
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_update_completed_
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_sample_start_
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_request/req
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_request/$entry
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_base_plus_offset/sum_rename_ack
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_base_plus_offset/sum_rename_req
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_base_plus_offset/$exit
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_base_plus_offset/$entry
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_final_index_sum_regn/ack
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_final_index_sum_regn/req
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_final_index_sum_regn/$exit
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_final_index_sum_regn/$entry
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_scale_0/scale_rename_ack
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_scale_0/scale_rename_req
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_scale_0/$exit
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_scale_0/$entry
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_resize_0/index_resize_ack
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_resize_0/index_resize_req
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_resize_0/$exit
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_resize_0/$entry
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_computed_0
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_scaled_0
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_index_resized_0
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_offset_calculated
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2380_Update/$exit
      -- CP-element group 693: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2384_root_address_calculated
      -- 
    ca_10701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 693_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2380_inst_ack_1, ack => minSumDecode_CP_6680_elements(693)); -- 
    req_10734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(693), ack => addr_of_2385_final_reg_req_0); -- 
    -- CP-element group 694:  transition  input  no-bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	693 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	704 
    -- CP-element group 694:  members (3) 
      -- CP-element group 694: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_request/ack
      -- CP-element group 694: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_request/$exit
      -- CP-element group 694: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_sample_completed_
      -- 
    ack_10735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2385_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(694)); -- 
    -- CP-element group 695:  transition  input  no-bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	691 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	704 
    -- CP-element group 695:  members (3) 
      -- CP-element group 695: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_complete/ack
      -- CP-element group 695: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_complete/$exit
      -- CP-element group 695: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2385_update_completed_
      -- 
    ack_10740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2385_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(695)); -- 
    -- CP-element group 696:  transition  input  no-bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	691 
    -- CP-element group 696: successors 
    -- CP-element group 696:  members (3) 
      -- CP-element group 696: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Sample/$exit
      -- CP-element group 696: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Sample/ra
      -- CP-element group 696: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_sample_completed_
      -- 
    ra_10749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 696_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_0, ack => minSumDecode_CP_6680_elements(696)); -- 
    -- CP-element group 697:  transition  input  output  no-bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	691 
    -- CP-element group 697: successors 
    -- CP-element group 697: 	702 
    -- CP-element group 697:  members (6) 
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_update_completed_
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Update/$exit
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/type_cast_2389_Update/ca
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_sample_start_
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Sample/$entry
      -- CP-element group 697: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Sample/rr
      -- 
    ca_10754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_1, ack => minSumDecode_CP_6680_elements(697)); -- 
    rr_10815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(697), ack => EQ_u32_u1_2404_inst_req_0); -- 
    -- CP-element group 698:  transition  input  no-bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	691 
    -- CP-element group 698: successors 
    -- CP-element group 698:  members (3) 
      -- CP-element group 698: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Sample/ra
      -- CP-element group 698: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Sample/$exit
      -- CP-element group 698: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_sample_completed_
      -- 
    ra_10763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2394_inst_ack_0, ack => minSumDecode_CP_6680_elements(698)); -- 
    -- CP-element group 699:  transition  input  output  no-bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	691 
    -- CP-element group 699: successors 
    -- CP-element group 699: 	700 
    -- CP-element group 699:  members (27) 
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Update/ca
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_Update/$exit
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_sample_start_
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/ADD_u64_u64_2394_update_completed_
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_root_address_calculated
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_offset_calculated
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_resized_0
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_scaled_0
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_computed_0
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_resize_0/$entry
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_resize_0/$exit
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_resize_0/index_resize_req
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_resize_0/index_resize_ack
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_scale_0/$entry
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_scale_0/$exit
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_scale_0/scale_rename_req
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_index_scale_0/scale_rename_ack
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_final_index_sum_regn/$entry
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_final_index_sum_regn/$exit
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_final_index_sum_regn/req
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_final_index_sum_regn/ack
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_base_plus_offset/$entry
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_base_plus_offset/$exit
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_base_plus_offset/sum_rename_req
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/array_obj_ref_2398_base_plus_offset/sum_rename_ack
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_request/$entry
      -- CP-element group 699: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_request/req
      -- 
    ca_10768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2394_inst_ack_1, ack => minSumDecode_CP_6680_elements(699)); -- 
    req_10801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(699), ack => addr_of_2399_final_reg_req_0); -- 
    -- CP-element group 700:  transition  input  no-bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	699 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	704 
    -- CP-element group 700:  members (3) 
      -- CP-element group 700: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_sample_completed_
      -- CP-element group 700: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_request/$exit
      -- CP-element group 700: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_request/ack
      -- 
    ack_10802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2399_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(700)); -- 
    -- CP-element group 701:  transition  input  no-bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	691 
    -- CP-element group 701: successors 
    -- CP-element group 701: 	704 
    -- CP-element group 701:  members (3) 
      -- CP-element group 701: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_update_completed_
      -- CP-element group 701: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_complete/$exit
      -- CP-element group 701: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/addr_of_2399_complete/ack
      -- 
    ack_10807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2399_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(701)); -- 
    -- CP-element group 702:  transition  input  no-bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	697 
    -- CP-element group 702: successors 
    -- CP-element group 702:  members (3) 
      -- CP-element group 702: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_sample_completed_
      -- CP-element group 702: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Sample/$exit
      -- CP-element group 702: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Sample/ra
      -- 
    ra_10816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2404_inst_ack_0, ack => minSumDecode_CP_6680_elements(702)); -- 
    -- CP-element group 703:  transition  input  no-bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	691 
    -- CP-element group 703: successors 
    -- CP-element group 703: 	704 
    -- CP-element group 703:  members (3) 
      -- CP-element group 703: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_update_completed_
      -- CP-element group 703: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Update/$exit
      -- CP-element group 703: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/EQ_u32_u1_2404_Update/ca
      -- 
    ca_10821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_2404_inst_ack_1, ack => minSumDecode_CP_6680_elements(703)); -- 
    -- CP-element group 704:  join  transition  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	694 
    -- CP-element group 704: 	695 
    -- CP-element group 704: 	700 
    -- CP-element group 704: 	701 
    -- CP-element group 704: 	703 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	80 
    -- CP-element group 704:  members (1) 
      -- CP-element group 704: 	 branch_block_stmt_1353/assign_stmt_2381_to_assign_stmt_2405/$exit
      -- 
    minSumDecode_cp_element_group_704: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_704"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(694) & minSumDecode_CP_6680_elements(695) & minSumDecode_CP_6680_elements(700) & minSumDecode_CP_6680_elements(701) & minSumDecode_CP_6680_elements(703);
      gj_minSumDecode_cp_element_group_704 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(704), clk => clk, reset => reset); --
    end block;
    -- CP-element group 705:  transition  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	80 
    -- CP-element group 705: successors 
    -- CP-element group 705:  members (1) 
      -- CP-element group 705: 	 branch_block_stmt_1353/if_stmt_2406_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(705) <= minSumDecode_CP_6680_elements(80);
    -- CP-element group 706:  transition  output  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	80 
    -- CP-element group 706: successors 
    -- CP-element group 706: 	707 
    -- CP-element group 706:  members (3) 
      -- CP-element group 706: 	 branch_block_stmt_1353/if_stmt_2406_eval_test/$entry
      -- CP-element group 706: 	 branch_block_stmt_1353/if_stmt_2406_eval_test/$exit
      -- CP-element group 706: 	 branch_block_stmt_1353/if_stmt_2406_eval_test/branch_req
      -- 
    branch_req_10829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(706), ack => if_stmt_2406_branch_req_0); -- 
    minSumDecode_CP_6680_elements(706) <= minSumDecode_CP_6680_elements(80);
    -- CP-element group 707:  branch  place  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	706 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	708 
    -- CP-element group 707: 	710 
    -- CP-element group 707:  members (1) 
      -- CP-element group 707: 	 branch_block_stmt_1353/R_iNsTr_140_2407_place
      -- 
    minSumDecode_CP_6680_elements(707) <= minSumDecode_CP_6680_elements(706);
    -- CP-element group 708:  transition  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	707 
    -- CP-element group 708: successors 
    -- CP-element group 708: 	709 
    -- CP-element group 708:  members (1) 
      -- CP-element group 708: 	 branch_block_stmt_1353/if_stmt_2406_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(708) <= minSumDecode_CP_6680_elements(707);
    -- CP-element group 709:  transition  input  no-bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	708 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	712 
    -- CP-element group 709:  members (2) 
      -- CP-element group 709: 	 branch_block_stmt_1353/if_stmt_2406_if_link/$exit
      -- CP-element group 709: 	 branch_block_stmt_1353/if_stmt_2406_if_link/if_choice_transition
      -- 
    if_choice_transition_10834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2406_branch_ack_1, ack => minSumDecode_CP_6680_elements(709)); -- 
    -- CP-element group 710:  transition  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	707 
    -- CP-element group 710: successors 
    -- CP-element group 710: 	711 
    -- CP-element group 710:  members (1) 
      -- CP-element group 710: 	 branch_block_stmt_1353/if_stmt_2406_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(710) <= minSumDecode_CP_6680_elements(707);
    -- CP-element group 711:  transition  input  no-bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	710 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	713 
    -- CP-element group 711:  members (2) 
      -- CP-element group 711: 	 branch_block_stmt_1353/if_stmt_2406_else_link/$exit
      -- CP-element group 711: 	 branch_block_stmt_1353/if_stmt_2406_else_link/else_choice_transition
      -- 
    else_choice_transition_10838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 711_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2406_branch_ack_0, ack => minSumDecode_CP_6680_elements(711)); -- 
    -- CP-element group 712:  place  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	709 
    -- CP-element group 712: successors 
    -- CP-element group 712: 	1124 
    -- CP-element group 712:  members (1) 
      -- CP-element group 712: 	 branch_block_stmt_1353/bb_41_bb_42
      -- 
    minSumDecode_CP_6680_elements(712) <= minSumDecode_CP_6680_elements(709);
    -- CP-element group 713:  place  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	711 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	1127 
    -- CP-element group 713:  members (1) 
      -- CP-element group 713: 	 branch_block_stmt_1353/bb_41_bb_43
      -- 
    minSumDecode_CP_6680_elements(713) <= minSumDecode_CP_6680_elements(711);
    -- CP-element group 714:  join  fork  transition  output  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	81 
    -- CP-element group 714: successors 
    -- CP-element group 714: 	715 
    -- CP-element group 714: 	716 
    -- CP-element group 714: 	718 
    -- CP-element group 714:  members (30) 
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_sample_start_
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_update_start_
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_address_calculated
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_word_address_calculated
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_root_address_calculated
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_address_resized
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_addr_resize/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_addr_resize/$exit
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_addr_resize/base_resize_req
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_addr_resize/base_resize_ack
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_plus_offset/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_plus_offset/$exit
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_plus_offset/sum_rename_req
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_base_plus_offset/sum_rename_ack
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_word_addrgen/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_word_addrgen/$exit
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_word_addrgen/root_register_req
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_word_addrgen/root_register_ack
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/word_0/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/word_0/rr
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/word_0/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/word_0/cr
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_update_start_
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Update/$entry
      -- CP-element group 714: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Update/cr
      -- 
    cr_10887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(714), ack => ptr_deref_2415_load_0_req_1); -- 
    rr_10876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(714), ack => ptr_deref_2415_load_0_req_0); -- 
    cr_10906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(714), ack => SUB_u16_u16_2420_inst_req_1); -- 
    minSumDecode_CP_6680_elements(714) <= minSumDecode_CP_6680_elements(81);
    -- CP-element group 715:  transition  input  no-bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	714 
    -- CP-element group 715: successors 
    -- CP-element group 715:  members (5) 
      -- CP-element group 715: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_sample_completed_
      -- CP-element group 715: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/$exit
      -- CP-element group 715: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/$exit
      -- CP-element group 715: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/word_0/$exit
      -- CP-element group 715: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Sample/word_access_start/word_0/ra
      -- 
    ra_10877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2415_load_0_ack_0, ack => minSumDecode_CP_6680_elements(715)); -- 
    -- CP-element group 716:  transition  input  output  no-bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	714 
    -- CP-element group 716: successors 
    -- CP-element group 716: 	717 
    -- CP-element group 716:  members (12) 
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_update_completed_
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/$exit
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/$exit
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/word_0/$exit
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/word_access_complete/word_0/ca
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/ptr_deref_2415_Merge/$entry
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/ptr_deref_2415_Merge/$exit
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/ptr_deref_2415_Merge/merge_req
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/ptr_deref_2415_Update/ptr_deref_2415_Merge/merge_ack
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_sample_start_
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Sample/$entry
      -- CP-element group 716: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Sample/rr
      -- 
    ca_10888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 716_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2415_load_0_ack_1, ack => minSumDecode_CP_6680_elements(716)); -- 
    rr_10901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(716), ack => SUB_u16_u16_2420_inst_req_0); -- 
    -- CP-element group 717:  transition  input  no-bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	716 
    -- CP-element group 717: successors 
    -- CP-element group 717:  members (3) 
      -- CP-element group 717: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_sample_completed_
      -- CP-element group 717: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Sample/$exit
      -- CP-element group 717: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Sample/ra
      -- 
    ra_10902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2420_inst_ack_0, ack => minSumDecode_CP_6680_elements(717)); -- 
    -- CP-element group 718:  transition  input  no-bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	714 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	82 
    -- CP-element group 718:  members (4) 
      -- CP-element group 718: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/$exit
      -- CP-element group 718: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_update_completed_
      -- CP-element group 718: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Update/$exit
      -- CP-element group 718: 	 branch_block_stmt_1353/assign_stmt_2416_to_assign_stmt_2421/SUB_u16_u16_2420_Update/ca
      -- 
    ca_10907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2420_inst_ack_1, ack => minSumDecode_CP_6680_elements(718)); -- 
    -- CP-element group 719:  join  fork  transition  output  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	83 
    -- CP-element group 719: successors 
    -- CP-element group 719: 	720 
    -- CP-element group 719: 	721 
    -- CP-element group 719: 	722 
    -- CP-element group 719: 	723 
    -- CP-element group 719: 	726 
    -- CP-element group 719:  members (56) 
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_sample_start_
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_update_start_
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_word_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_root_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_address_resized
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_addr_resize/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_addr_resize/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_addr_resize/base_resize_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_addr_resize/base_resize_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_plus_offset/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_plus_offset/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_plus_offset/sum_rename_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_base_plus_offset/sum_rename_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_word_addrgen/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_word_addrgen/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_word_addrgen/root_register_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_word_addrgen/root_register_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/word_0/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/word_0/rr
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/word_0/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/word_0/cr
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_sample_start_
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_update_start_
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_word_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_root_address_calculated
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_address_resized
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_addr_resize/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_addr_resize/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_addr_resize/base_resize_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_addr_resize/base_resize_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_plus_offset/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_plus_offset/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_plus_offset/sum_rename_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_base_plus_offset/sum_rename_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_word_addrgen/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_word_addrgen/$exit
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_word_addrgen/root_register_req
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_word_addrgen/root_register_ack
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/word_0/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/word_0/rr
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/word_0/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/word_0/cr
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_update_start_
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Update/$entry
      -- CP-element group 719: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Update/cr
      -- 
    cr_10954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(719), ack => ptr_deref_2426_load_0_req_1); -- 
    rr_10943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(719), ack => ptr_deref_2426_load_0_req_0); -- 
    cr_11004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(719), ack => ptr_deref_2430_load_0_req_1); -- 
    rr_10993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(719), ack => ptr_deref_2430_load_0_req_0); -- 
    cr_11023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(719), ack => SUB_u16_u16_2435_inst_req_1); -- 
    minSumDecode_CP_6680_elements(719) <= minSumDecode_CP_6680_elements(83);
    -- CP-element group 720:  transition  input  no-bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	719 
    -- CP-element group 720: successors 
    -- CP-element group 720:  members (5) 
      -- CP-element group 720: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_sample_completed_
      -- CP-element group 720: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/$exit
      -- CP-element group 720: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/$exit
      -- CP-element group 720: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/word_0/$exit
      -- CP-element group 720: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Sample/word_access_start/word_0/ra
      -- 
    ra_10944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 720_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2426_load_0_ack_0, ack => minSumDecode_CP_6680_elements(720)); -- 
    -- CP-element group 721:  transition  input  no-bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	719 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	724 
    -- CP-element group 721:  members (9) 
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_update_completed_
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/$exit
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/$exit
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/word_0/$exit
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/word_access_complete/word_0/ca
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/ptr_deref_2426_Merge/$entry
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/ptr_deref_2426_Merge/$exit
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/ptr_deref_2426_Merge/merge_req
      -- CP-element group 721: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2426_Update/ptr_deref_2426_Merge/merge_ack
      -- 
    ca_10955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 721_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2426_load_0_ack_1, ack => minSumDecode_CP_6680_elements(721)); -- 
    -- CP-element group 722:  transition  input  no-bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	719 
    -- CP-element group 722: successors 
    -- CP-element group 722:  members (5) 
      -- CP-element group 722: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_sample_completed_
      -- CP-element group 722: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/$exit
      -- CP-element group 722: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/$exit
      -- CP-element group 722: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/word_0/$exit
      -- CP-element group 722: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Sample/word_access_start/word_0/ra
      -- 
    ra_10994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2430_load_0_ack_0, ack => minSumDecode_CP_6680_elements(722)); -- 
    -- CP-element group 723:  transition  input  no-bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	719 
    -- CP-element group 723: successors 
    -- CP-element group 723: 	724 
    -- CP-element group 723:  members (9) 
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_update_completed_
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/$exit
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/$exit
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/word_0/$exit
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/word_access_complete/word_0/ca
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/ptr_deref_2430_Merge/$entry
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/ptr_deref_2430_Merge/$exit
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/ptr_deref_2430_Merge/merge_req
      -- CP-element group 723: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/ptr_deref_2430_Update/ptr_deref_2430_Merge/merge_ack
      -- 
    ca_11005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 723_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2430_load_0_ack_1, ack => minSumDecode_CP_6680_elements(723)); -- 
    -- CP-element group 724:  join  transition  output  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	721 
    -- CP-element group 724: 	723 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	725 
    -- CP-element group 724:  members (3) 
      -- CP-element group 724: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_sample_start_
      -- CP-element group 724: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Sample/$entry
      -- CP-element group 724: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Sample/rr
      -- 
    rr_11018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(724), ack => SUB_u16_u16_2435_inst_req_0); -- 
    minSumDecode_cp_element_group_724: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_724"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(721) & minSumDecode_CP_6680_elements(723);
      gj_minSumDecode_cp_element_group_724 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(724), clk => clk, reset => reset); --
    end block;
    -- CP-element group 725:  transition  input  no-bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	724 
    -- CP-element group 725: successors 
    -- CP-element group 725:  members (3) 
      -- CP-element group 725: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_sample_completed_
      -- CP-element group 725: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Sample/$exit
      -- CP-element group 725: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Sample/ra
      -- 
    ra_11019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2435_inst_ack_0, ack => minSumDecode_CP_6680_elements(725)); -- 
    -- CP-element group 726:  transition  input  no-bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	719 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	84 
    -- CP-element group 726:  members (4) 
      -- CP-element group 726: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/$exit
      -- CP-element group 726: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_update_completed_
      -- CP-element group 726: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Update/$exit
      -- CP-element group 726: 	 branch_block_stmt_1353/assign_stmt_2427_to_assign_stmt_2436/SUB_u16_u16_2435_Update/ca
      -- 
    ca_11024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 726_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2435_inst_ack_1, ack => minSumDecode_CP_6680_elements(726)); -- 
    -- CP-element group 727:  fork  transition  output  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	85 
    -- CP-element group 727: successors 
    -- CP-element group 727: 	728 
    -- CP-element group 727: 	729 
    -- CP-element group 727:  members (7) 
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/$entry
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_sample_start_
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_update_start_
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Sample/$entry
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Sample/rr
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Update/$entry
      -- CP-element group 727: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Update/cr
      -- 
    rr_11035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(727), ack => EQ_u16_u1_2456_inst_req_0); -- 
    cr_11040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(727), ack => EQ_u16_u1_2456_inst_req_1); -- 
    minSumDecode_CP_6680_elements(727) <= minSumDecode_CP_6680_elements(85);
    -- CP-element group 728:  transition  input  no-bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	727 
    -- CP-element group 728: successors 
    -- CP-element group 728:  members (3) 
      -- CP-element group 728: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_sample_completed_
      -- CP-element group 728: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Sample/$exit
      -- CP-element group 728: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Sample/ra
      -- 
    ra_11036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2456_inst_ack_0, ack => minSumDecode_CP_6680_elements(728)); -- 
    -- CP-element group 729:  transition  input  no-bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	727 
    -- CP-element group 729: successors 
    -- CP-element group 729: 	86 
    -- CP-element group 729:  members (4) 
      -- CP-element group 729: 	 branch_block_stmt_1353/assign_stmt_2457/$exit
      -- CP-element group 729: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_update_completed_
      -- CP-element group 729: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Update/$exit
      -- CP-element group 729: 	 branch_block_stmt_1353/assign_stmt_2457/EQ_u16_u1_2456_Update/ca
      -- 
    ca_11041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 729_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2456_inst_ack_1, ack => minSumDecode_CP_6680_elements(729)); -- 
    -- CP-element group 730:  transition  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	86 
    -- CP-element group 730: successors 
    -- CP-element group 730:  members (1) 
      -- CP-element group 730: 	 branch_block_stmt_1353/if_stmt_2458_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(730) <= minSumDecode_CP_6680_elements(86);
    -- CP-element group 731:  transition  output  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	86 
    -- CP-element group 731: successors 
    -- CP-element group 731: 	732 
    -- CP-element group 731:  members (3) 
      -- CP-element group 731: 	 branch_block_stmt_1353/if_stmt_2458_eval_test/$entry
      -- CP-element group 731: 	 branch_block_stmt_1353/if_stmt_2458_eval_test/$exit
      -- CP-element group 731: 	 branch_block_stmt_1353/if_stmt_2458_eval_test/branch_req
      -- 
    branch_req_11049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(731), ack => if_stmt_2458_branch_req_0); -- 
    minSumDecode_CP_6680_elements(731) <= minSumDecode_CP_6680_elements(86);
    -- CP-element group 732:  branch  place  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	731 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732: 	735 
    -- CP-element group 732:  members (1) 
      -- CP-element group 732: 	 branch_block_stmt_1353/R_iNsTr_150_2459_place
      -- 
    minSumDecode_CP_6680_elements(732) <= minSumDecode_CP_6680_elements(731);
    -- CP-element group 733:  transition  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733: 	734 
    -- CP-element group 733:  members (1) 
      -- CP-element group 733: 	 branch_block_stmt_1353/if_stmt_2458_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(733) <= minSumDecode_CP_6680_elements(732);
    -- CP-element group 734:  transition  input  no-bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	733 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	737 
    -- CP-element group 734:  members (2) 
      -- CP-element group 734: 	 branch_block_stmt_1353/if_stmt_2458_if_link/$exit
      -- CP-element group 734: 	 branch_block_stmt_1353/if_stmt_2458_if_link/if_choice_transition
      -- 
    if_choice_transition_11054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2458_branch_ack_1, ack => minSumDecode_CP_6680_elements(734)); -- 
    -- CP-element group 735:  transition  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	732 
    -- CP-element group 735: successors 
    -- CP-element group 735: 	736 
    -- CP-element group 735:  members (1) 
      -- CP-element group 735: 	 branch_block_stmt_1353/if_stmt_2458_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(735) <= minSumDecode_CP_6680_elements(732);
    -- CP-element group 736:  transition  input  no-bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	735 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	738 
    -- CP-element group 736:  members (2) 
      -- CP-element group 736: 	 branch_block_stmt_1353/if_stmt_2458_else_link/$exit
      -- CP-element group 736: 	 branch_block_stmt_1353/if_stmt_2458_else_link/else_choice_transition
      -- 
    else_choice_transition_11058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 736_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2458_branch_ack_0, ack => minSumDecode_CP_6680_elements(736)); -- 
    -- CP-element group 737:  place  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	734 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	1167 
    -- CP-element group 737:  members (1) 
      -- CP-element group 737: 	 branch_block_stmt_1353/bb_44_xx_x_crit_edgex_xi
      -- 
    minSumDecode_CP_6680_elements(737) <= minSumDecode_CP_6680_elements(734);
    -- CP-element group 738:  place  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	736 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	1151 
    -- CP-element group 738:  members (1) 
      -- CP-element group 738: 	 branch_block_stmt_1353/bb_44_bbx_xnphx_xi36
      -- 
    minSumDecode_CP_6680_elements(738) <= minSumDecode_CP_6680_elements(736);
    -- CP-element group 739:  fork  transition  output  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	87 
    -- CP-element group 739: successors 
    -- CP-element group 739: 	740 
    -- CP-element group 739: 	741 
    -- CP-element group 739:  members (7) 
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/$entry
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_sample_start_
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_update_start_
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Sample/$entry
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Sample/rr
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Update/cr
      -- 
    rr_11071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(739), ack => ADD_u16_u16_2469_inst_req_0); -- 
    cr_11076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(739), ack => ADD_u16_u16_2469_inst_req_1); -- 
    minSumDecode_CP_6680_elements(739) <= minSumDecode_CP_6680_elements(87);
    -- CP-element group 740:  transition  input  no-bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	739 
    -- CP-element group 740: successors 
    -- CP-element group 740:  members (3) 
      -- CP-element group 740: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_sample_completed_
      -- CP-element group 740: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Sample/$exit
      -- CP-element group 740: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Sample/ra
      -- 
    ra_11072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2469_inst_ack_0, ack => minSumDecode_CP_6680_elements(740)); -- 
    -- CP-element group 741:  transition  input  no-bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	739 
    -- CP-element group 741: successors 
    -- CP-element group 741: 	88 
    -- CP-element group 741:  members (4) 
      -- CP-element group 741: 	 branch_block_stmt_1353/assign_stmt_2470/$exit
      -- CP-element group 741: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_update_completed_
      -- CP-element group 741: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Update/$exit
      -- CP-element group 741: 	 branch_block_stmt_1353/assign_stmt_2470/ADD_u16_u16_2469_Update/ca
      -- 
    ca_11077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 741_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2469_inst_ack_1, ack => minSumDecode_CP_6680_elements(741)); -- 
    -- CP-element group 742:  fork  transition  output  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	89 
    -- CP-element group 742: successors 
    -- CP-element group 742: 	743 
    -- CP-element group 742: 	744 
    -- CP-element group 742: 	746 
    -- CP-element group 742: 	748 
    -- CP-element group 742: 	750 
    -- CP-element group 742: 	752 
    -- CP-element group 742: 	754 
    -- CP-element group 742: 	756 
    -- CP-element group 742: 	758 
    -- CP-element group 742: 	760 
    -- CP-element group 742: 	762 
    -- CP-element group 742: 	764 
    -- CP-element group 742: 	767 
    -- CP-element group 742: 	769 
    -- CP-element group 742: 	772 
    -- CP-element group 742: 	773 
    -- CP-element group 742: 	774 
    -- CP-element group 742: 	776 
    -- CP-element group 742:  members (63) 
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_sample_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Sample/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Sample/rr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_complete/req
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/word_0/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/word_0/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_complete/req
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/word_0/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/word_0/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_complete/req
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/word_0/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/word_0/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_complete/req
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/word_0/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/word_0/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_sample_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Sample/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Sample/rr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Update/cr
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_update_start_
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Update/$entry
      -- CP-element group 742: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Update/cr
      -- 
    rr_11088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u16_u16_2484_inst_req_0); -- 
    cr_11093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u16_u16_2484_inst_req_1); -- 
    cr_11107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => type_cast_2488_inst_req_1); -- 
    cr_11121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u64_u64_2494_inst_req_1); -- 
    req_11160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => addr_of_2499_final_reg_req_1); -- 
    cr_11205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ptr_deref_2503_load_0_req_1); -- 
    cr_11224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u16_u16_2509_inst_req_1); -- 
    cr_11238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => type_cast_2513_inst_req_1); -- 
    req_11277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => addr_of_2518_final_reg_req_1); -- 
    cr_11322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ptr_deref_2522_load_0_req_1); -- 
    req_11366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => addr_of_2527_final_reg_req_1); -- 
    cr_11411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ptr_deref_2531_load_0_req_1); -- 
    cr_11430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => SUB_f32_f32_2536_inst_req_1); -- 
    req_11469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => addr_of_2541_final_reg_req_1); -- 
    cr_11519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ptr_deref_2544_store_0_req_1); -- 
    rr_11528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u16_u16_2551_inst_req_0); -- 
    cr_11533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => ADD_u16_u16_2551_inst_req_1); -- 
    cr_11547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(742), ack => EQ_u16_u1_2556_inst_req_1); -- 
    minSumDecode_CP_6680_elements(742) <= minSumDecode_CP_6680_elements(89);
    -- CP-element group 743:  transition  input  no-bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	742 
    -- CP-element group 743: successors 
    -- CP-element group 743:  members (3) 
      -- CP-element group 743: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_sample_completed_
      -- CP-element group 743: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Sample/$exit
      -- CP-element group 743: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Sample/ra
      -- 
    ra_11089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 743_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2484_inst_ack_0, ack => minSumDecode_CP_6680_elements(743)); -- 
    -- CP-element group 744:  transition  input  output  no-bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	742 
    -- CP-element group 744: successors 
    -- CP-element group 744: 	745 
    -- CP-element group 744:  members (6) 
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_update_completed_
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Update/$exit
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2484_Update/ca
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_sample_start_
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Sample/$entry
      -- CP-element group 744: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Sample/rr
      -- 
    ca_11094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 744_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2484_inst_ack_1, ack => minSumDecode_CP_6680_elements(744)); -- 
    rr_11102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(744), ack => type_cast_2488_inst_req_0); -- 
    -- CP-element group 745:  transition  input  no-bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	744 
    -- CP-element group 745: successors 
    -- CP-element group 745:  members (3) 
      -- CP-element group 745: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_sample_completed_
      -- CP-element group 745: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Sample/$exit
      -- CP-element group 745: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Sample/ra
      -- 
    ra_11103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 745_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2488_inst_ack_0, ack => minSumDecode_CP_6680_elements(745)); -- 
    -- CP-element group 746:  fork  transition  input  output  no-bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	742 
    -- CP-element group 746: successors 
    -- CP-element group 746: 	747 
    -- CP-element group 746: 	761 
    -- CP-element group 746: 	768 
    -- CP-element group 746:  members (54) 
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_update_completed_
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Update/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2488_Update/ca
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_sample_start_
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Sample/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Sample/rr
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_sample_start_
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_root_address_calculated
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_offset_calculated
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_resized_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_scaled_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_computed_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_resize_0/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_resize_0/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_resize_0/index_resize_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_resize_0/index_resize_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_scale_0/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_scale_0/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_scale_0/scale_rename_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_index_scale_0/scale_rename_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_final_index_sum_regn/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_final_index_sum_regn/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_final_index_sum_regn/req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_final_index_sum_regn/ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_base_plus_offset/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_base_plus_offset/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_base_plus_offset/sum_rename_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2526_base_plus_offset/sum_rename_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_request/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_request/req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_sample_start_
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_root_address_calculated
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_offset_calculated
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_resized_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_scaled_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_computed_0
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_resize_0/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_resize_0/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_resize_0/index_resize_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_resize_0/index_resize_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_scale_0/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_scale_0/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_scale_0/scale_rename_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_index_scale_0/scale_rename_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_final_index_sum_regn/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_final_index_sum_regn/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_final_index_sum_regn/req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_final_index_sum_regn/ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_base_plus_offset/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_base_plus_offset/$exit
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_base_plus_offset/sum_rename_req
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2540_base_plus_offset/sum_rename_ack
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_request/$entry
      -- CP-element group 746: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_request/req
      -- 
    ca_11108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 746_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2488_inst_ack_1, ack => minSumDecode_CP_6680_elements(746)); -- 
    rr_11116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(746), ack => ADD_u64_u64_2494_inst_req_0); -- 
    req_11361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(746), ack => addr_of_2527_final_reg_req_0); -- 
    req_11464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(746), ack => addr_of_2541_final_reg_req_0); -- 
    -- CP-element group 747:  transition  input  no-bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	746 
    -- CP-element group 747: successors 
    -- CP-element group 747:  members (3) 
      -- CP-element group 747: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_sample_completed_
      -- CP-element group 747: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Sample/$exit
      -- CP-element group 747: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Sample/ra
      -- 
    ra_11117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2494_inst_ack_0, ack => minSumDecode_CP_6680_elements(747)); -- 
    -- CP-element group 748:  transition  input  output  no-bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	742 
    -- CP-element group 748: successors 
    -- CP-element group 748: 	749 
    -- CP-element group 748:  members (27) 
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_update_completed_
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Update/$exit
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u64_u64_2494_Update/ca
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_sample_start_
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_root_address_calculated
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_offset_calculated
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_resized_0
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_scaled_0
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_computed_0
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_resize_0/$entry
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_resize_0/$exit
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_resize_0/index_resize_req
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_resize_0/index_resize_ack
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_scale_0/$entry
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_scale_0/$exit
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_scale_0/scale_rename_req
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_index_scale_0/scale_rename_ack
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_final_index_sum_regn/$entry
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_final_index_sum_regn/$exit
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_final_index_sum_regn/req
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_final_index_sum_regn/ack
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_base_plus_offset/$entry
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_base_plus_offset/$exit
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_base_plus_offset/sum_rename_req
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2498_base_plus_offset/sum_rename_ack
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_request/$entry
      -- CP-element group 748: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_request/req
      -- 
    ca_11122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2494_inst_ack_1, ack => minSumDecode_CP_6680_elements(748)); -- 
    req_11155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(748), ack => addr_of_2499_final_reg_req_0); -- 
    -- CP-element group 749:  transition  input  no-bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	748 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	777 
    -- CP-element group 749:  members (3) 
      -- CP-element group 749: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_sample_completed_
      -- CP-element group 749: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_request/$exit
      -- CP-element group 749: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_request/ack
      -- 
    ack_11156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 749_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2499_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(749)); -- 
    -- CP-element group 750:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	742 
    -- CP-element group 750: successors 
    -- CP-element group 750: 	751 
    -- CP-element group 750:  members (24) 
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_update_completed_
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_complete/$exit
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2499_complete/ack
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_sample_start_
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_address_calculated
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_word_address_calculated
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_root_address_calculated
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_address_resized
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_addr_resize/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_addr_resize/$exit
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_addr_resize/base_resize_req
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_addr_resize/base_resize_ack
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_plus_offset/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_plus_offset/$exit
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_plus_offset/sum_rename_req
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_base_plus_offset/sum_rename_ack
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_word_addrgen/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_word_addrgen/$exit
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_word_addrgen/root_register_req
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_word_addrgen/root_register_ack
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/word_0/$entry
      -- CP-element group 750: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/word_0/rr
      -- 
    ack_11161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2499_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(750)); -- 
    rr_11194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(750), ack => ptr_deref_2503_load_0_req_0); -- 
    -- CP-element group 751:  transition  input  no-bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	750 
    -- CP-element group 751: successors 
    -- CP-element group 751:  members (5) 
      -- CP-element group 751: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_sample_completed_
      -- CP-element group 751: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/$exit
      -- CP-element group 751: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/$exit
      -- CP-element group 751: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/word_0/$exit
      -- CP-element group 751: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Sample/word_access_start/word_0/ra
      -- 
    ra_11195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2503_load_0_ack_0, ack => minSumDecode_CP_6680_elements(751)); -- 
    -- CP-element group 752:  transition  input  output  no-bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	742 
    -- CP-element group 752: successors 
    -- CP-element group 752: 	753 
    -- CP-element group 752:  members (12) 
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_update_completed_
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/$exit
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/$exit
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/word_0/$exit
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/word_access_complete/word_0/ca
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/ptr_deref_2503_Merge/$entry
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/ptr_deref_2503_Merge/$exit
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/ptr_deref_2503_Merge/merge_req
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2503_Update/ptr_deref_2503_Merge/merge_ack
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_sample_start_
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Sample/$entry
      -- CP-element group 752: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Sample/rr
      -- 
    ca_11206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 752_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2503_load_0_ack_1, ack => minSumDecode_CP_6680_elements(752)); -- 
    rr_11219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(752), ack => ADD_u16_u16_2509_inst_req_0); -- 
    -- CP-element group 753:  transition  input  no-bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	752 
    -- CP-element group 753: successors 
    -- CP-element group 753:  members (3) 
      -- CP-element group 753: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_sample_completed_
      -- CP-element group 753: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Sample/$exit
      -- CP-element group 753: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Sample/ra
      -- 
    ra_11220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 753_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2509_inst_ack_0, ack => minSumDecode_CP_6680_elements(753)); -- 
    -- CP-element group 754:  transition  input  output  no-bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	742 
    -- CP-element group 754: successors 
    -- CP-element group 754: 	755 
    -- CP-element group 754:  members (6) 
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_update_completed_
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Update/$exit
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2509_Update/ca
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_sample_start_
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Sample/$entry
      -- CP-element group 754: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Sample/rr
      -- 
    ca_11225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2509_inst_ack_1, ack => minSumDecode_CP_6680_elements(754)); -- 
    rr_11233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(754), ack => type_cast_2513_inst_req_0); -- 
    -- CP-element group 755:  transition  input  no-bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	754 
    -- CP-element group 755: successors 
    -- CP-element group 755:  members (3) 
      -- CP-element group 755: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_sample_completed_
      -- CP-element group 755: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Sample/$exit
      -- CP-element group 755: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Sample/ra
      -- 
    ra_11234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 755_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_0, ack => minSumDecode_CP_6680_elements(755)); -- 
    -- CP-element group 756:  transition  input  output  no-bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	742 
    -- CP-element group 756: successors 
    -- CP-element group 756: 	757 
    -- CP-element group 756:  members (27) 
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_scaled_0
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_update_completed_
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Update/$exit
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/type_cast_2513_Update/ca
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_sample_start_
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_root_address_calculated
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_offset_calculated
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_resized_0
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_computed_0
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_resize_0/$entry
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_resize_0/$exit
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_resize_0/index_resize_req
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_resize_0/index_resize_ack
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_scale_0/$entry
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_scale_0/$exit
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_scale_0/scale_rename_req
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_index_scale_0/scale_rename_ack
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_final_index_sum_regn/$entry
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_final_index_sum_regn/$exit
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_final_index_sum_regn/req
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_final_index_sum_regn/ack
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_base_plus_offset/$entry
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_base_plus_offset/$exit
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_base_plus_offset/sum_rename_req
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/array_obj_ref_2517_base_plus_offset/sum_rename_ack
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_request/$entry
      -- CP-element group 756: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_request/req
      -- 
    ca_11239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 756_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_1, ack => minSumDecode_CP_6680_elements(756)); -- 
    req_11272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(756), ack => addr_of_2518_final_reg_req_0); -- 
    -- CP-element group 757:  transition  input  no-bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	756 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	777 
    -- CP-element group 757:  members (3) 
      -- CP-element group 757: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_sample_completed_
      -- CP-element group 757: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_request/$exit
      -- CP-element group 757: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_request/ack
      -- 
    ack_11273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2518_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(757)); -- 
    -- CP-element group 758:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	742 
    -- CP-element group 758: successors 
    -- CP-element group 758: 	759 
    -- CP-element group 758:  members (24) 
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_update_completed_
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_complete/$exit
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2518_complete/ack
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_sample_start_
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_address_calculated
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_word_address_calculated
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_root_address_calculated
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_address_resized
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_addr_resize/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_addr_resize/$exit
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_addr_resize/base_resize_req
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_addr_resize/base_resize_ack
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_plus_offset/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_plus_offset/$exit
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_plus_offset/sum_rename_req
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_base_plus_offset/sum_rename_ack
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_word_addrgen/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_word_addrgen/$exit
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_word_addrgen/root_register_req
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_word_addrgen/root_register_ack
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/word_0/$entry
      -- CP-element group 758: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/word_0/rr
      -- 
    ack_11278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2518_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(758)); -- 
    rr_11311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(758), ack => ptr_deref_2522_load_0_req_0); -- 
    -- CP-element group 759:  transition  input  no-bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	758 
    -- CP-element group 759: successors 
    -- CP-element group 759:  members (5) 
      -- CP-element group 759: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_sample_completed_
      -- CP-element group 759: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/$exit
      -- CP-element group 759: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/$exit
      -- CP-element group 759: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/word_0/$exit
      -- CP-element group 759: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Sample/word_access_start/word_0/ra
      -- 
    ra_11312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 759_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2522_load_0_ack_0, ack => minSumDecode_CP_6680_elements(759)); -- 
    -- CP-element group 760:  transition  input  no-bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	742 
    -- CP-element group 760: successors 
    -- CP-element group 760: 	765 
    -- CP-element group 760:  members (9) 
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_update_completed_
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/$exit
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/$exit
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/word_0/$exit
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/word_access_complete/word_0/ca
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/ptr_deref_2522_Merge/$entry
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/ptr_deref_2522_Merge/$exit
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/ptr_deref_2522_Merge/merge_req
      -- CP-element group 760: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2522_Update/ptr_deref_2522_Merge/merge_ack
      -- 
    ca_11323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2522_load_0_ack_1, ack => minSumDecode_CP_6680_elements(760)); -- 
    -- CP-element group 761:  transition  input  no-bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	746 
    -- CP-element group 761: successors 
    -- CP-element group 761: 	777 
    -- CP-element group 761:  members (3) 
      -- CP-element group 761: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_sample_completed_
      -- CP-element group 761: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_request/$exit
      -- CP-element group 761: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_request/ack
      -- 
    ack_11362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2527_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(761)); -- 
    -- CP-element group 762:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	742 
    -- CP-element group 762: successors 
    -- CP-element group 762: 	763 
    -- CP-element group 762:  members (24) 
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_update_completed_
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_complete/$exit
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2527_complete/ack
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_sample_start_
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_address_calculated
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_word_address_calculated
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_root_address_calculated
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_address_resized
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_addr_resize/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_addr_resize/$exit
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_addr_resize/base_resize_req
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_addr_resize/base_resize_ack
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_plus_offset/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_plus_offset/$exit
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_plus_offset/sum_rename_req
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_base_plus_offset/sum_rename_ack
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_word_addrgen/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_word_addrgen/$exit
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_word_addrgen/root_register_req
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_word_addrgen/root_register_ack
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/word_0/$entry
      -- CP-element group 762: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/word_0/rr
      -- 
    ack_11367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 762_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2527_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(762)); -- 
    rr_11400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(762), ack => ptr_deref_2531_load_0_req_0); -- 
    -- CP-element group 763:  transition  input  no-bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	762 
    -- CP-element group 763: successors 
    -- CP-element group 763:  members (5) 
      -- CP-element group 763: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_sample_completed_
      -- CP-element group 763: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/$exit
      -- CP-element group 763: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/$exit
      -- CP-element group 763: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/word_0/$exit
      -- CP-element group 763: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Sample/word_access_start/word_0/ra
      -- 
    ra_11401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 763_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2531_load_0_ack_0, ack => minSumDecode_CP_6680_elements(763)); -- 
    -- CP-element group 764:  transition  input  no-bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	742 
    -- CP-element group 764: successors 
    -- CP-element group 764: 	765 
    -- CP-element group 764:  members (9) 
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_update_completed_
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/$exit
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/$exit
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/word_0/$exit
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/word_access_complete/word_0/ca
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/ptr_deref_2531_Merge/$entry
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/ptr_deref_2531_Merge/$exit
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/ptr_deref_2531_Merge/merge_req
      -- CP-element group 764: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2531_Update/ptr_deref_2531_Merge/merge_ack
      -- 
    ca_11412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 764_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2531_load_0_ack_1, ack => minSumDecode_CP_6680_elements(764)); -- 
    -- CP-element group 765:  join  transition  output  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	760 
    -- CP-element group 765: 	764 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	766 
    -- CP-element group 765:  members (3) 
      -- CP-element group 765: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_sample_start_
      -- CP-element group 765: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Sample/$entry
      -- CP-element group 765: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Sample/rr
      -- 
    rr_11425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(765), ack => SUB_f32_f32_2536_inst_req_0); -- 
    minSumDecode_cp_element_group_765: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_765"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(760) & minSumDecode_CP_6680_elements(764);
      gj_minSumDecode_cp_element_group_765 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(765), clk => clk, reset => reset); --
    end block;
    -- CP-element group 766:  transition  input  no-bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	765 
    -- CP-element group 766: successors 
    -- CP-element group 766:  members (3) 
      -- CP-element group 766: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_sample_completed_
      -- CP-element group 766: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Sample/$exit
      -- CP-element group 766: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Sample/ra
      -- 
    ra_11426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 766_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2536_inst_ack_0, ack => minSumDecode_CP_6680_elements(766)); -- 
    -- CP-element group 767:  transition  input  no-bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	742 
    -- CP-element group 767: successors 
    -- CP-element group 767: 	770 
    -- CP-element group 767:  members (3) 
      -- CP-element group 767: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_update_completed_
      -- CP-element group 767: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Update/$exit
      -- CP-element group 767: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/SUB_f32_f32_2536_Update/ca
      -- 
    ca_11431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_f32_f32_2536_inst_ack_1, ack => minSumDecode_CP_6680_elements(767)); -- 
    -- CP-element group 768:  transition  input  no-bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	746 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	777 
    -- CP-element group 768:  members (3) 
      -- CP-element group 768: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_sample_completed_
      -- CP-element group 768: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_request/$exit
      -- CP-element group 768: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_request/ack
      -- 
    ack_11465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 768_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2541_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(768)); -- 
    -- CP-element group 769:  fork  transition  input  no-bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	742 
    -- CP-element group 769: successors 
    -- CP-element group 769: 	770 
    -- CP-element group 769:  members (19) 
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_update_completed_
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_complete/$exit
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/addr_of_2541_complete/ack
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_address_calculated
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_word_address_calculated
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_root_address_calculated
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_address_resized
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_addr_resize/$entry
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_addr_resize/$exit
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_addr_resize/base_resize_req
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_addr_resize/base_resize_ack
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_plus_offset/$entry
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_plus_offset/$exit
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_plus_offset/sum_rename_req
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_base_plus_offset/sum_rename_ack
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_word_addrgen/$entry
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_word_addrgen/$exit
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_word_addrgen/root_register_req
      -- CP-element group 769: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_word_addrgen/root_register_ack
      -- 
    ack_11470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 769_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2541_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(769)); -- 
    -- CP-element group 770:  join  transition  output  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	767 
    -- CP-element group 770: 	769 
    -- CP-element group 770: successors 
    -- CP-element group 770: 	771 
    -- CP-element group 770:  members (9) 
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_sample_start_
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/$entry
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/ptr_deref_2544_Split/$entry
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/ptr_deref_2544_Split/$exit
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/ptr_deref_2544_Split/split_req
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/ptr_deref_2544_Split/split_ack
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/$entry
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/word_0/$entry
      -- CP-element group 770: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/word_0/rr
      -- 
    rr_11508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(770), ack => ptr_deref_2544_store_0_req_0); -- 
    minSumDecode_cp_element_group_770: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_770"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(767) & minSumDecode_CP_6680_elements(769);
      gj_minSumDecode_cp_element_group_770 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(770), clk => clk, reset => reset); --
    end block;
    -- CP-element group 771:  transition  input  no-bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	770 
    -- CP-element group 771: successors 
    -- CP-element group 771:  members (5) 
      -- CP-element group 771: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_sample_completed_
      -- CP-element group 771: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/$exit
      -- CP-element group 771: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/$exit
      -- CP-element group 771: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/word_0/$exit
      -- CP-element group 771: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Sample/word_access_start/word_0/ra
      -- 
    ra_11509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 771_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2544_store_0_ack_0, ack => minSumDecode_CP_6680_elements(771)); -- 
    -- CP-element group 772:  transition  input  no-bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	742 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	777 
    -- CP-element group 772:  members (5) 
      -- CP-element group 772: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_update_completed_
      -- CP-element group 772: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/$exit
      -- CP-element group 772: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/$exit
      -- CP-element group 772: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/word_0/$exit
      -- CP-element group 772: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ptr_deref_2544_Update/word_access_complete/word_0/ca
      -- 
    ca_11520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 772_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2544_store_0_ack_1, ack => minSumDecode_CP_6680_elements(772)); -- 
    -- CP-element group 773:  transition  input  no-bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	742 
    -- CP-element group 773: successors 
    -- CP-element group 773:  members (3) 
      -- CP-element group 773: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_sample_completed_
      -- CP-element group 773: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Sample/$exit
      -- CP-element group 773: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Sample/ra
      -- 
    ra_11529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 773_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2551_inst_ack_0, ack => minSumDecode_CP_6680_elements(773)); -- 
    -- CP-element group 774:  transition  input  output  no-bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	742 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	775 
    -- CP-element group 774:  members (6) 
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_update_completed_
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Update/$exit
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/ADD_u16_u16_2551_Update/ca
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_sample_start_
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Sample/$entry
      -- CP-element group 774: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Sample/rr
      -- 
    ca_11534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 774_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2551_inst_ack_1, ack => minSumDecode_CP_6680_elements(774)); -- 
    rr_11542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(774), ack => EQ_u16_u1_2556_inst_req_0); -- 
    -- CP-element group 775:  transition  input  no-bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	774 
    -- CP-element group 775: successors 
    -- CP-element group 775:  members (3) 
      -- CP-element group 775: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_sample_completed_
      -- CP-element group 775: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Sample/$exit
      -- CP-element group 775: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Sample/ra
      -- 
    ra_11543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 775_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2556_inst_ack_0, ack => minSumDecode_CP_6680_elements(775)); -- 
    -- CP-element group 776:  transition  input  no-bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	742 
    -- CP-element group 776: successors 
    -- CP-element group 776: 	777 
    -- CP-element group 776:  members (3) 
      -- CP-element group 776: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_update_completed_
      -- CP-element group 776: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Update/$exit
      -- CP-element group 776: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/EQ_u16_u1_2556_Update/ca
      -- 
    ca_11548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 776_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2556_inst_ack_1, ack => minSumDecode_CP_6680_elements(776)); -- 
    -- CP-element group 777:  join  transition  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	749 
    -- CP-element group 777: 	757 
    -- CP-element group 777: 	761 
    -- CP-element group 777: 	768 
    -- CP-element group 777: 	772 
    -- CP-element group 777: 	776 
    -- CP-element group 777: successors 
    -- CP-element group 777: 	90 
    -- CP-element group 777:  members (1) 
      -- CP-element group 777: 	 branch_block_stmt_1353/assign_stmt_2485_to_assign_stmt_2557/$exit
      -- 
    minSumDecode_cp_element_group_777: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_777"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(749) & minSumDecode_CP_6680_elements(757) & minSumDecode_CP_6680_elements(761) & minSumDecode_CP_6680_elements(768) & minSumDecode_CP_6680_elements(772) & minSumDecode_CP_6680_elements(776);
      gj_minSumDecode_cp_element_group_777 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(777), clk => clk, reset => reset); --
    end block;
    -- CP-element group 778:  transition  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	90 
    -- CP-element group 778: successors 
    -- CP-element group 778:  members (1) 
      -- CP-element group 778: 	 branch_block_stmt_1353/if_stmt_2558_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(778) <= minSumDecode_CP_6680_elements(90);
    -- CP-element group 779:  transition  output  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	90 
    -- CP-element group 779: successors 
    -- CP-element group 779: 	780 
    -- CP-element group 779:  members (3) 
      -- CP-element group 779: 	 branch_block_stmt_1353/if_stmt_2558_eval_test/$entry
      -- CP-element group 779: 	 branch_block_stmt_1353/if_stmt_2558_eval_test/$exit
      -- CP-element group 779: 	 branch_block_stmt_1353/if_stmt_2558_eval_test/branch_req
      -- 
    branch_req_11556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(779), ack => if_stmt_2558_branch_req_0); -- 
    minSumDecode_CP_6680_elements(779) <= minSumDecode_CP_6680_elements(90);
    -- CP-element group 780:  branch  place  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	779 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	781 
    -- CP-element group 780: 	783 
    -- CP-element group 780:  members (1) 
      -- CP-element group 780: 	 branch_block_stmt_1353/R_exitcond5_2559_place
      -- 
    minSumDecode_CP_6680_elements(780) <= minSumDecode_CP_6680_elements(779);
    -- CP-element group 781:  transition  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	780 
    -- CP-element group 781: successors 
    -- CP-element group 781: 	782 
    -- CP-element group 781:  members (1) 
      -- CP-element group 781: 	 branch_block_stmt_1353/if_stmt_2558_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(781) <= minSumDecode_CP_6680_elements(780);
    -- CP-element group 782:  transition  input  no-bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	781 
    -- CP-element group 782: successors 
    -- CP-element group 782: 	785 
    -- CP-element group 782:  members (2) 
      -- CP-element group 782: 	 branch_block_stmt_1353/if_stmt_2558_if_link/$exit
      -- CP-element group 782: 	 branch_block_stmt_1353/if_stmt_2558_if_link/if_choice_transition
      -- 
    if_choice_transition_11561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 782_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2558_branch_ack_1, ack => minSumDecode_CP_6680_elements(782)); -- 
    -- CP-element group 783:  transition  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	780 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	784 
    -- CP-element group 783:  members (1) 
      -- CP-element group 783: 	 branch_block_stmt_1353/if_stmt_2558_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(783) <= minSumDecode_CP_6680_elements(780);
    -- CP-element group 784:  transition  input  no-bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	783 
    -- CP-element group 784: successors 
    -- CP-element group 784: 	786 
    -- CP-element group 784:  members (2) 
      -- CP-element group 784: 	 branch_block_stmt_1353/if_stmt_2558_else_link/$exit
      -- CP-element group 784: 	 branch_block_stmt_1353/if_stmt_2558_else_link/else_choice_transition
      -- 
    else_choice_transition_11565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 784_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2558_branch_ack_0, ack => minSumDecode_CP_6680_elements(784)); -- 
    -- CP-element group 785:  place  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	782 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	1164 
    -- CP-element group 785:  members (1) 
      -- CP-element group 785: 	 branch_block_stmt_1353/bb_46_xx_x_crit_edgex_xix_xloopexit
      -- 
    minSumDecode_CP_6680_elements(785) <= minSumDecode_CP_6680_elements(782);
    -- CP-element group 786:  place  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	784 
    -- CP-element group 786: successors 
    -- CP-element group 786: 	1154 
    -- CP-element group 786:  members (1) 
      -- CP-element group 786: 	 branch_block_stmt_1353/bb_46_bb_46
      -- 
    minSumDecode_CP_6680_elements(786) <= minSumDecode_CP_6680_elements(784);
    -- CP-element group 787:  fork  transition  output  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	92 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	788 
    -- CP-element group 787: 	789 
    -- CP-element group 787: 	791 
    -- CP-element group 787:  members (10) 
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/$entry
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_sample_start_
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_update_start_
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Sample/$entry
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Sample/rr
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Update/$entry
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Update/cr
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_update_start_
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Update/$entry
      -- CP-element group 787: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Update/cr
      -- 
    rr_11578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(787), ack => ADD_u64_u64_2571_inst_req_0); -- 
    cr_11583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(787), ack => ADD_u64_u64_2571_inst_req_1); -- 
    cr_11597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(787), ack => EQ_u64_u1_2576_inst_req_1); -- 
    minSumDecode_CP_6680_elements(787) <= minSumDecode_CP_6680_elements(92);
    -- CP-element group 788:  transition  input  no-bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	787 
    -- CP-element group 788: successors 
    -- CP-element group 788:  members (3) 
      -- CP-element group 788: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_sample_completed_
      -- CP-element group 788: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Sample/$exit
      -- CP-element group 788: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Sample/ra
      -- 
    ra_11579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 788_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2571_inst_ack_0, ack => minSumDecode_CP_6680_elements(788)); -- 
    -- CP-element group 789:  transition  input  output  no-bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	787 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	790 
    -- CP-element group 789:  members (6) 
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_update_completed_
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Update/$exit
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/ADD_u64_u64_2571_Update/ca
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_sample_start_
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Sample/$entry
      -- CP-element group 789: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Sample/rr
      -- 
    ca_11584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 789_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2571_inst_ack_1, ack => minSumDecode_CP_6680_elements(789)); -- 
    rr_11592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(789), ack => EQ_u64_u1_2576_inst_req_0); -- 
    -- CP-element group 790:  transition  input  no-bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	789 
    -- CP-element group 790: successors 
    -- CP-element group 790:  members (3) 
      -- CP-element group 790: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_sample_completed_
      -- CP-element group 790: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Sample/$exit
      -- CP-element group 790: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Sample/ra
      -- 
    ra_11593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 790_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2576_inst_ack_0, ack => minSumDecode_CP_6680_elements(790)); -- 
    -- CP-element group 791:  transition  input  no-bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	787 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	93 
    -- CP-element group 791:  members (4) 
      -- CP-element group 791: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/$exit
      -- CP-element group 791: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_update_completed_
      -- CP-element group 791: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Update/$exit
      -- CP-element group 791: 	 branch_block_stmt_1353/assign_stmt_2572_to_assign_stmt_2577/EQ_u64_u1_2576_Update/ca
      -- 
    ca_11598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 791_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u64_u1_2576_inst_ack_1, ack => minSumDecode_CP_6680_elements(791)); -- 
    -- CP-element group 792:  transition  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	93 
    -- CP-element group 792: successors 
    -- CP-element group 792:  members (1) 
      -- CP-element group 792: 	 branch_block_stmt_1353/if_stmt_2578_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(792) <= minSumDecode_CP_6680_elements(93);
    -- CP-element group 793:  transition  output  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	93 
    -- CP-element group 793: successors 
    -- CP-element group 793: 	794 
    -- CP-element group 793:  members (3) 
      -- CP-element group 793: 	 branch_block_stmt_1353/if_stmt_2578_eval_test/$entry
      -- CP-element group 793: 	 branch_block_stmt_1353/if_stmt_2578_eval_test/$exit
      -- CP-element group 793: 	 branch_block_stmt_1353/if_stmt_2578_eval_test/branch_req
      -- 
    branch_req_11606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(793), ack => if_stmt_2578_branch_req_0); -- 
    minSumDecode_CP_6680_elements(793) <= minSumDecode_CP_6680_elements(93);
    -- CP-element group 794:  branch  place  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	793 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	795 
    -- CP-element group 794: 	797 
    -- CP-element group 794:  members (1) 
      -- CP-element group 794: 	 branch_block_stmt_1353/R_exitcond6_2579_place
      -- 
    minSumDecode_CP_6680_elements(794) <= minSumDecode_CP_6680_elements(793);
    -- CP-element group 795:  transition  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	794 
    -- CP-element group 795: successors 
    -- CP-element group 795: 	796 
    -- CP-element group 795:  members (1) 
      -- CP-element group 795: 	 branch_block_stmt_1353/if_stmt_2578_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(795) <= minSumDecode_CP_6680_elements(794);
    -- CP-element group 796:  transition  input  no-bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	795 
    -- CP-element group 796: successors 
    -- CP-element group 796: 	799 
    -- CP-element group 796:  members (2) 
      -- CP-element group 796: 	 branch_block_stmt_1353/if_stmt_2578_if_link/$exit
      -- CP-element group 796: 	 branch_block_stmt_1353/if_stmt_2578_if_link/if_choice_transition
      -- 
    if_choice_transition_11611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 796_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2578_branch_ack_1, ack => minSumDecode_CP_6680_elements(796)); -- 
    -- CP-element group 797:  transition  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	794 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	798 
    -- CP-element group 797:  members (1) 
      -- CP-element group 797: 	 branch_block_stmt_1353/if_stmt_2578_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(797) <= minSumDecode_CP_6680_elements(794);
    -- CP-element group 798:  transition  input  no-bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	797 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	800 
    -- CP-element group 798:  members (2) 
      -- CP-element group 798: 	 branch_block_stmt_1353/if_stmt_2578_else_link/$exit
      -- CP-element group 798: 	 branch_block_stmt_1353/if_stmt_2578_else_link/else_choice_transition
      -- 
    else_choice_transition_11615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 798_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2578_branch_ack_0, ack => minSumDecode_CP_6680_elements(798)); -- 
    -- CP-element group 799:  place  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	796 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	1171 
    -- CP-element group 799:  members (1) 
      -- CP-element group 799: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_updateMessagex_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(799) <= minSumDecode_CP_6680_elements(796);
    -- CP-element group 800:  place  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	798 
    -- CP-element group 800: successors 
    -- CP-element group 800: 	1117 
    -- CP-element group 800:  members (1) 
      -- CP-element group 800: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41
      -- 
    minSumDecode_CP_6680_elements(800) <= minSumDecode_CP_6680_elements(798);
    -- CP-element group 801:  fork  transition  output  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	95 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	802 
    -- CP-element group 801: 	803 
    -- CP-element group 801:  members (7) 
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/$entry
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_sample_start_
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_update_start_
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Sample/$entry
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Sample/rr
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Update/$entry
      -- CP-element group 801: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Update/cr
      -- 
    rr_11628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(801), ack => ADD_u16_u16_2591_inst_req_0); -- 
    cr_11633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(801), ack => ADD_u16_u16_2591_inst_req_1); -- 
    minSumDecode_CP_6680_elements(801) <= minSumDecode_CP_6680_elements(95);
    -- CP-element group 802:  transition  input  no-bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	801 
    -- CP-element group 802: successors 
    -- CP-element group 802:  members (3) 
      -- CP-element group 802: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_sample_completed_
      -- CP-element group 802: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Sample/$exit
      -- CP-element group 802: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Sample/ra
      -- 
    ra_11629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 802_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2591_inst_ack_0, ack => minSumDecode_CP_6680_elements(802)); -- 
    -- CP-element group 803:  transition  input  no-bypass 
    -- CP-element group 803: predecessors 
    -- CP-element group 803: 	801 
    -- CP-element group 803: successors 
    -- CP-element group 803: 	96 
    -- CP-element group 803:  members (4) 
      -- CP-element group 803: 	 branch_block_stmt_1353/assign_stmt_2592/$exit
      -- CP-element group 803: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_update_completed_
      -- CP-element group 803: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Update/$exit
      -- CP-element group 803: 	 branch_block_stmt_1353/assign_stmt_2592/ADD_u16_u16_2591_Update/ca
      -- 
    ca_11634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 803_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_2591_inst_ack_1, ack => minSumDecode_CP_6680_elements(803)); -- 
    -- CP-element group 804:  fork  transition  output  bypass 
    -- CP-element group 804: predecessors 
    -- CP-element group 804: 	97 
    -- CP-element group 804: successors 
    -- CP-element group 804: 	805 
    -- CP-element group 804: 	806 
    -- CP-element group 804: 	807 
    -- CP-element group 804: 	808 
    -- CP-element group 804:  members (23) 
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_sample_start_
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_update_start_
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_word_address_calculated
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_root_address_calculated
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/STORE_Nitr_required_2608_Split/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/STORE_Nitr_required_2608_Split/$exit
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/STORE_Nitr_required_2608_Split/split_req
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/STORE_Nitr_required_2608_Split/split_ack
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/word_0/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/word_0/rr
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/word_0/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/word_0/cr
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_sample_start_
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_update_start_
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Sample/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Sample/rr
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Update/$entry
      -- CP-element group 804: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Update/cr
      -- 
    cr_11669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(804), ack => STORE_Nitr_required_2608_store_0_req_1); -- 
    rr_11658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(804), ack => STORE_Nitr_required_2608_store_0_req_0); -- 
    rr_11678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(804), ack => EQ_u16_u1_2615_inst_req_0); -- 
    cr_11683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(804), ack => EQ_u16_u1_2615_inst_req_1); -- 
    minSumDecode_CP_6680_elements(804) <= minSumDecode_CP_6680_elements(97);
    -- CP-element group 805:  transition  input  no-bypass 
    -- CP-element group 805: predecessors 
    -- CP-element group 805: 	804 
    -- CP-element group 805: successors 
    -- CP-element group 805:  members (5) 
      -- CP-element group 805: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_sample_completed_
      -- CP-element group 805: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/$exit
      -- CP-element group 805: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/$exit
      -- CP-element group 805: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/word_0/$exit
      -- CP-element group 805: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Sample/word_access_start/word_0/ra
      -- 
    ra_11659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 805_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_Nitr_required_2608_store_0_ack_0, ack => minSumDecode_CP_6680_elements(805)); -- 
    -- CP-element group 806:  transition  input  no-bypass 
    -- CP-element group 806: predecessors 
    -- CP-element group 806: 	804 
    -- CP-element group 806: successors 
    -- CP-element group 806: 	809 
    -- CP-element group 806:  members (5) 
      -- CP-element group 806: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_update_completed_
      -- CP-element group 806: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/$exit
      -- CP-element group 806: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/$exit
      -- CP-element group 806: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/word_0/$exit
      -- CP-element group 806: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/STORE_Nitr_required_2608_Update/word_access_complete/word_0/ca
      -- 
    ca_11670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 806_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_Nitr_required_2608_store_0_ack_1, ack => minSumDecode_CP_6680_elements(806)); -- 
    -- CP-element group 807:  transition  input  no-bypass 
    -- CP-element group 807: predecessors 
    -- CP-element group 807: 	804 
    -- CP-element group 807: successors 
    -- CP-element group 807:  members (3) 
      -- CP-element group 807: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_sample_completed_
      -- CP-element group 807: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Sample/$exit
      -- CP-element group 807: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Sample/ra
      -- 
    ra_11679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 807_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2615_inst_ack_0, ack => minSumDecode_CP_6680_elements(807)); -- 
    -- CP-element group 808:  transition  input  no-bypass 
    -- CP-element group 808: predecessors 
    -- CP-element group 808: 	804 
    -- CP-element group 808: successors 
    -- CP-element group 808: 	809 
    -- CP-element group 808:  members (3) 
      -- CP-element group 808: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_update_completed_
      -- CP-element group 808: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Update/$exit
      -- CP-element group 808: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/EQ_u16_u1_2615_Update/ca
      -- 
    ca_11684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 808_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u16_u1_2615_inst_ack_1, ack => minSumDecode_CP_6680_elements(808)); -- 
    -- CP-element group 809:  join  transition  bypass 
    -- CP-element group 809: predecessors 
    -- CP-element group 809: 	806 
    -- CP-element group 809: 	808 
    -- CP-element group 809: successors 
    -- CP-element group 809: 	98 
    -- CP-element group 809:  members (1) 
      -- CP-element group 809: 	 branch_block_stmt_1353/assign_stmt_2610_to_assign_stmt_2616/$exit
      -- 
    minSumDecode_cp_element_group_809: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_809"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(806) & minSumDecode_CP_6680_elements(808);
      gj_minSumDecode_cp_element_group_809 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(809), clk => clk, reset => reset); --
    end block;
    -- CP-element group 810:  transition  bypass 
    -- CP-element group 810: predecessors 
    -- CP-element group 810: 	98 
    -- CP-element group 810: successors 
    -- CP-element group 810:  members (1) 
      -- CP-element group 810: 	 branch_block_stmt_1353/if_stmt_2617_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(810) <= minSumDecode_CP_6680_elements(98);
    -- CP-element group 811:  transition  output  bypass 
    -- CP-element group 811: predecessors 
    -- CP-element group 811: 	98 
    -- CP-element group 811: successors 
    -- CP-element group 811: 	812 
    -- CP-element group 811:  members (3) 
      -- CP-element group 811: 	 branch_block_stmt_1353/if_stmt_2617_eval_test/$entry
      -- CP-element group 811: 	 branch_block_stmt_1353/if_stmt_2617_eval_test/$exit
      -- CP-element group 811: 	 branch_block_stmt_1353/if_stmt_2617_eval_test/branch_req
      -- 
    branch_req_11692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(811), ack => if_stmt_2617_branch_req_0); -- 
    minSumDecode_CP_6680_elements(811) <= minSumDecode_CP_6680_elements(98);
    -- CP-element group 812:  branch  place  bypass 
    -- CP-element group 812: predecessors 
    -- CP-element group 812: 	811 
    -- CP-element group 812: successors 
    -- CP-element group 812: 	813 
    -- CP-element group 812: 	815 
    -- CP-element group 812:  members (1) 
      -- CP-element group 812: 	 branch_block_stmt_1353/R_iNsTr_43_2618_place
      -- 
    minSumDecode_CP_6680_elements(812) <= minSumDecode_CP_6680_elements(811);
    -- CP-element group 813:  transition  bypass 
    -- CP-element group 813: predecessors 
    -- CP-element group 813: 	812 
    -- CP-element group 813: successors 
    -- CP-element group 813: 	814 
    -- CP-element group 813:  members (1) 
      -- CP-element group 813: 	 branch_block_stmt_1353/if_stmt_2617_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(813) <= minSumDecode_CP_6680_elements(812);
    -- CP-element group 814:  transition  input  no-bypass 
    -- CP-element group 814: predecessors 
    -- CP-element group 814: 	813 
    -- CP-element group 814: successors 
    -- CP-element group 814: 	817 
    -- CP-element group 814:  members (2) 
      -- CP-element group 814: 	 branch_block_stmt_1353/if_stmt_2617_if_link/$exit
      -- CP-element group 814: 	 branch_block_stmt_1353/if_stmt_2617_if_link/if_choice_transition
      -- 
    if_choice_transition_11697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 814_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2617_branch_ack_1, ack => minSumDecode_CP_6680_elements(814)); -- 
    -- CP-element group 815:  transition  bypass 
    -- CP-element group 815: predecessors 
    -- CP-element group 815: 	812 
    -- CP-element group 815: successors 
    -- CP-element group 815: 	816 
    -- CP-element group 815:  members (1) 
      -- CP-element group 815: 	 branch_block_stmt_1353/if_stmt_2617_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(815) <= minSumDecode_CP_6680_elements(812);
    -- CP-element group 816:  transition  input  no-bypass 
    -- CP-element group 816: predecessors 
    -- CP-element group 816: 	815 
    -- CP-element group 816: successors 
    -- CP-element group 816: 	818 
    -- CP-element group 816:  members (2) 
      -- CP-element group 816: 	 branch_block_stmt_1353/if_stmt_2617_else_link/$exit
      -- CP-element group 816: 	 branch_block_stmt_1353/if_stmt_2617_else_link/else_choice_transition
      -- 
    else_choice_transition_11701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 816_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2617_branch_ack_0, ack => minSumDecode_CP_6680_elements(816)); -- 
    -- CP-element group 817:  place  bypass 
    -- CP-element group 817: predecessors 
    -- CP-element group 817: 	814 
    -- CP-element group 817: successors 
    -- CP-element group 817: 	1215 
    -- CP-element group 817:  members (1) 
      -- CP-element group 817: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit
      -- 
    minSumDecode_CP_6680_elements(817) <= minSumDecode_CP_6680_elements(814);
    -- CP-element group 818:  place  bypass 
    -- CP-element group 818: predecessors 
    -- CP-element group 818: 	816 
    -- CP-element group 818: successors 
    -- CP-element group 818: 	1199 
    -- CP-element group 818:  members (1) 
      -- CP-element group 818: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_bbx_xnphx_xi13x_xpreheader
      -- 
    minSumDecode_CP_6680_elements(818) <= minSumDecode_CP_6680_elements(816);
    -- CP-element group 819:  fork  transition  output  bypass 
    -- CP-element group 819: predecessors 
    -- CP-element group 819: 	100 
    -- CP-element group 819: successors 
    -- CP-element group 819: 	820 
    -- CP-element group 819: 	821 
    -- CP-element group 819: 	822 
    -- CP-element group 819: 	823 
    -- CP-element group 819: 	825 
    -- CP-element group 819: 	826 
    -- CP-element group 819: 	827 
    -- CP-element group 819: 	829 
    -- CP-element group 819:  members (48) 
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_sample_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_update_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_root_address_calculated
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_offset_calculated
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_resized_0
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_scaled_0
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_computed_0
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_resize_0/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_resize_0/$exit
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_resize_0/index_resize_req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_resize_0/index_resize_ack
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_scale_0/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_scale_0/$exit
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_scale_0/scale_rename_req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_index_scale_0/scale_rename_ack
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn/$exit
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn/req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn/ack
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/$exit
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/sum_rename_req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/sum_rename_ack
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_request/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_request/req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_complete/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_complete/req
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_sample_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_update_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Sample/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Sample/rr
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Update/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Update/cr
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_update_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Update/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Update/cr
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_sample_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_update_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Sample/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Sample/rr
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Update/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Update/cr
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_update_start_
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/word_0/$entry
      -- CP-element group 819: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/word_0/cr
      -- 
    req_11744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => addr_of_2637_final_reg_req_1); -- 
    req_11739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => addr_of_2637_final_reg_req_0); -- 
    rr_11753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => ADD_u64_u64_2643_inst_req_0); -- 
    cr_11758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => ADD_u64_u64_2643_inst_req_1); -- 
    cr_11772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => type_cast_2647_inst_req_1); -- 
    rr_11781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => ADD_u64_u64_2653_inst_req_0); -- 
    cr_11786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => ADD_u64_u64_2653_inst_req_1); -- 
    cr_11831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(819), ack => ptr_deref_2657_load_0_req_1); -- 
    minSumDecode_CP_6680_elements(819) <= minSumDecode_CP_6680_elements(100);
    -- CP-element group 820:  transition  input  no-bypass 
    -- CP-element group 820: predecessors 
    -- CP-element group 820: 	819 
    -- CP-element group 820: successors 
    -- CP-element group 820: 	830 
    -- CP-element group 820:  members (3) 
      -- CP-element group 820: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_sample_completed_
      -- CP-element group 820: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_request/$exit
      -- CP-element group 820: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_request/ack
      -- 
    ack_11740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 820_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2637_final_reg_ack_0, ack => minSumDecode_CP_6680_elements(820)); -- 
    -- CP-element group 821:  join  fork  transition  input  output  no-bypass 
    -- CP-element group 821: predecessors 
    -- CP-element group 821: 	819 
    -- CP-element group 821: successors 
    -- CP-element group 821: 	828 
    -- CP-element group 821:  members (24) 
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_update_completed_
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_complete/$exit
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/addr_of_2637_complete/ack
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_sample_start_
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_address_calculated
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_word_address_calculated
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_root_address_calculated
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_address_resized
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_addr_resize/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_addr_resize/$exit
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_addr_resize/base_resize_req
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_addr_resize/base_resize_ack
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_plus_offset/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_plus_offset/$exit
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_plus_offset/sum_rename_req
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_base_plus_offset/sum_rename_ack
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_word_addrgen/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_word_addrgen/$exit
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_word_addrgen/root_register_req
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_word_addrgen/root_register_ack
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/word_0/$entry
      -- CP-element group 821: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/word_0/rr
      -- 
    ack_11745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 821_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2637_final_reg_ack_1, ack => minSumDecode_CP_6680_elements(821)); -- 
    rr_11820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(821), ack => ptr_deref_2657_load_0_req_0); -- 
    -- CP-element group 822:  transition  input  no-bypass 
    -- CP-element group 822: predecessors 
    -- CP-element group 822: 	819 
    -- CP-element group 822: successors 
    -- CP-element group 822:  members (3) 
      -- CP-element group 822: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_sample_completed_
      -- CP-element group 822: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Sample/$exit
      -- CP-element group 822: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Sample/ra
      -- 
    ra_11754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 822_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2643_inst_ack_0, ack => minSumDecode_CP_6680_elements(822)); -- 
    -- CP-element group 823:  transition  input  output  no-bypass 
    -- CP-element group 823: predecessors 
    -- CP-element group 823: 	819 
    -- CP-element group 823: successors 
    -- CP-element group 823: 	824 
    -- CP-element group 823:  members (6) 
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_update_completed_
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Update/$exit
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2643_Update/ca
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_sample_start_
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Sample/$entry
      -- CP-element group 823: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Sample/rr
      -- 
    ca_11759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 823_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2643_inst_ack_1, ack => minSumDecode_CP_6680_elements(823)); -- 
    rr_11767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(823), ack => type_cast_2647_inst_req_0); -- 
    -- CP-element group 824:  transition  input  no-bypass 
    -- CP-element group 824: predecessors 
    -- CP-element group 824: 	823 
    -- CP-element group 824: successors 
    -- CP-element group 824:  members (3) 
      -- CP-element group 824: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_sample_completed_
      -- CP-element group 824: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Sample/$exit
      -- CP-element group 824: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Sample/ra
      -- 
    ra_11768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 824_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_0, ack => minSumDecode_CP_6680_elements(824)); -- 
    -- CP-element group 825:  transition  input  no-bypass 
    -- CP-element group 825: predecessors 
    -- CP-element group 825: 	819 
    -- CP-element group 825: successors 
    -- CP-element group 825: 	830 
    -- CP-element group 825:  members (3) 
      -- CP-element group 825: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_update_completed_
      -- CP-element group 825: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Update/$exit
      -- CP-element group 825: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/type_cast_2647_Update/ca
      -- 
    ca_11773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 825_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_1, ack => minSumDecode_CP_6680_elements(825)); -- 
    -- CP-element group 826:  transition  input  no-bypass 
    -- CP-element group 826: predecessors 
    -- CP-element group 826: 	819 
    -- CP-element group 826: successors 
    -- CP-element group 826:  members (3) 
      -- CP-element group 826: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_sample_completed_
      -- CP-element group 826: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Sample/$exit
      -- CP-element group 826: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Sample/ra
      -- 
    ra_11782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 826_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2653_inst_ack_0, ack => minSumDecode_CP_6680_elements(826)); -- 
    -- CP-element group 827:  transition  input  no-bypass 
    -- CP-element group 827: predecessors 
    -- CP-element group 827: 	819 
    -- CP-element group 827: successors 
    -- CP-element group 827: 	830 
    -- CP-element group 827:  members (3) 
      -- CP-element group 827: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_update_completed_
      -- CP-element group 827: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Update/$exit
      -- CP-element group 827: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ADD_u64_u64_2653_Update/ca
      -- 
    ca_11787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 827_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2653_inst_ack_1, ack => minSumDecode_CP_6680_elements(827)); -- 
    -- CP-element group 828:  transition  input  no-bypass 
    -- CP-element group 828: predecessors 
    -- CP-element group 828: 	821 
    -- CP-element group 828: successors 
    -- CP-element group 828:  members (5) 
      -- CP-element group 828: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_sample_completed_
      -- CP-element group 828: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/$exit
      -- CP-element group 828: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/$exit
      -- CP-element group 828: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/word_0/$exit
      -- CP-element group 828: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Sample/word_access_start/word_0/ra
      -- 
    ra_11821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 828_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2657_load_0_ack_0, ack => minSumDecode_CP_6680_elements(828)); -- 
    -- CP-element group 829:  transition  input  no-bypass 
    -- CP-element group 829: predecessors 
    -- CP-element group 829: 	819 
    -- CP-element group 829: successors 
    -- CP-element group 829: 	830 
    -- CP-element group 829:  members (9) 
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_update_completed_
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/$exit
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/$exit
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/word_0/$exit
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/word_access_complete/word_0/ca
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/ptr_deref_2657_Merge/$entry
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/ptr_deref_2657_Merge/$exit
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/ptr_deref_2657_Merge/merge_req
      -- CP-element group 829: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/ptr_deref_2657_Update/ptr_deref_2657_Merge/merge_ack
      -- 
    ca_11832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 829_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2657_load_0_ack_1, ack => minSumDecode_CP_6680_elements(829)); -- 
    -- CP-element group 830:  join  transition  bypass 
    -- CP-element group 830: predecessors 
    -- CP-element group 830: 	820 
    -- CP-element group 830: 	825 
    -- CP-element group 830: 	827 
    -- CP-element group 830: 	829 
    -- CP-element group 830: successors 
    -- CP-element group 830: 	101 
    -- CP-element group 830:  members (1) 
      -- CP-element group 830: 	 branch_block_stmt_1353/assign_stmt_2638_to_assign_stmt_2658/$exit
      -- 
    minSumDecode_cp_element_group_830: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_830"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(820) & minSumDecode_CP_6680_elements(825) & minSumDecode_CP_6680_elements(827) & minSumDecode_CP_6680_elements(829);
      gj_minSumDecode_cp_element_group_830 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(830), clk => clk, reset => reset); --
    end block;
    -- CP-element group 831:  transition  output  bypass 
    -- CP-element group 831: predecessors 
    -- CP-element group 831: 	101 
    -- CP-element group 831: successors 
    -- CP-element group 831: 	832 
    -- CP-element group 831:  members (4) 
      -- CP-element group 831: 	 branch_block_stmt_1353/assign_stmt_2661/$entry
      -- CP-element group 831: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_sample_start_
      -- CP-element group 831: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Sample/$entry
      -- CP-element group 831: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Sample/req
      -- 
    req_11848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(831), ack => WPIPE_code_block_decoded_2659_inst_req_0); -- 
    minSumDecode_CP_6680_elements(831) <= minSumDecode_CP_6680_elements(101);
    -- CP-element group 832:  transition  input  output  no-bypass 
    -- CP-element group 832: predecessors 
    -- CP-element group 832: 	831 
    -- CP-element group 832: successors 
    -- CP-element group 832: 	833 
    -- CP-element group 832:  members (6) 
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_sample_completed_
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_update_start_
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Sample/$exit
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Sample/ack
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Update/$entry
      -- CP-element group 832: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Update/req
      -- 
    ack_11849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 832_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_code_block_decoded_2659_inst_ack_0, ack => minSumDecode_CP_6680_elements(832)); -- 
    req_11853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(832), ack => WPIPE_code_block_decoded_2659_inst_req_1); -- 
    -- CP-element group 833:  transition  input  no-bypass 
    -- CP-element group 833: predecessors 
    -- CP-element group 833: 	832 
    -- CP-element group 833: successors 
    -- CP-element group 833: 	102 
    -- CP-element group 833:  members (4) 
      -- CP-element group 833: 	 branch_block_stmt_1353/assign_stmt_2661/$exit
      -- CP-element group 833: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_update_completed_
      -- CP-element group 833: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Update/$exit
      -- CP-element group 833: 	 branch_block_stmt_1353/assign_stmt_2661/WPIPE_code_block_decoded_2659_Update/ack
      -- 
    ack_11854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 833_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_code_block_decoded_2659_inst_ack_1, ack => minSumDecode_CP_6680_elements(833)); -- 
    -- CP-element group 834:  fork  transition  output  bypass 
    -- CP-element group 834: predecessors 
    -- CP-element group 834: 	102 
    -- CP-element group 834: successors 
    -- CP-element group 834: 	835 
    -- CP-element group 834: 	836 
    -- CP-element group 834: 	838 
    -- CP-element group 834: 	840 
    -- CP-element group 834:  members (19) 
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_sample_start_
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_update_start_
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_word_address_calculated
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_root_address_calculated
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/word_0/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/word_0/rr
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/word_0/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/word_0/cr
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_update_start_
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Update/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Update/cr
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_update_start_
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Update/$entry
      -- CP-element group 834: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Update/cr
      -- 
    cr_11884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(834), ack => LOAD_ncols_2663_load_0_req_1); -- 
    rr_11873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(834), ack => LOAD_ncols_2663_load_0_req_0); -- 
    cr_11903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(834), ack => type_cast_2667_inst_req_1); -- 
    cr_11917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(834), ack => SLT_i32_u1_2675_inst_req_1); -- 
    minSumDecode_CP_6680_elements(834) <= minSumDecode_CP_6680_elements(102);
    -- CP-element group 835:  transition  input  no-bypass 
    -- CP-element group 835: predecessors 
    -- CP-element group 835: 	834 
    -- CP-element group 835: successors 
    -- CP-element group 835:  members (5) 
      -- CP-element group 835: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_sample_completed_
      -- CP-element group 835: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/$exit
      -- CP-element group 835: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/$exit
      -- CP-element group 835: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/word_0/$exit
      -- CP-element group 835: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Sample/word_access_start/word_0/ra
      -- 
    ra_11874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 835_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_2663_load_0_ack_0, ack => minSumDecode_CP_6680_elements(835)); -- 
    -- CP-element group 836:  transition  input  output  no-bypass 
    -- CP-element group 836: predecessors 
    -- CP-element group 836: 	834 
    -- CP-element group 836: successors 
    -- CP-element group 836: 	837 
    -- CP-element group 836:  members (12) 
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_update_completed_
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/$exit
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/$exit
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/word_0/$exit
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/word_access_complete/word_0/ca
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/LOAD_ncols_2663_Merge/$entry
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/LOAD_ncols_2663_Merge/$exit
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/LOAD_ncols_2663_Merge/merge_req
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/LOAD_ncols_2663_Update/LOAD_ncols_2663_Merge/merge_ack
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_sample_start_
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Sample/$entry
      -- CP-element group 836: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Sample/rr
      -- 
    ca_11885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 836_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ncols_2663_load_0_ack_1, ack => minSumDecode_CP_6680_elements(836)); -- 
    rr_11898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(836), ack => type_cast_2667_inst_req_0); -- 
    -- CP-element group 837:  transition  input  no-bypass 
    -- CP-element group 837: predecessors 
    -- CP-element group 837: 	836 
    -- CP-element group 837: successors 
    -- CP-element group 837:  members (3) 
      -- CP-element group 837: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_sample_completed_
      -- CP-element group 837: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Sample/$exit
      -- CP-element group 837: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Sample/ra
      -- 
    ra_11899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 837_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_0, ack => minSumDecode_CP_6680_elements(837)); -- 
    -- CP-element group 838:  transition  input  output  no-bypass 
    -- CP-element group 838: predecessors 
    -- CP-element group 838: 	834 
    -- CP-element group 838: successors 
    -- CP-element group 838: 	839 
    -- CP-element group 838:  members (6) 
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_update_completed_
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Update/$exit
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/type_cast_2667_Update/ca
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_sample_start_
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Sample/$entry
      -- CP-element group 838: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Sample/rr
      -- 
    ca_11904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 838_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_1, ack => minSumDecode_CP_6680_elements(838)); -- 
    rr_11912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(838), ack => SLT_i32_u1_2675_inst_req_0); -- 
    -- CP-element group 839:  transition  input  no-bypass 
    -- CP-element group 839: predecessors 
    -- CP-element group 839: 	838 
    -- CP-element group 839: successors 
    -- CP-element group 839:  members (3) 
      -- CP-element group 839: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_sample_completed_
      -- CP-element group 839: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Sample/$exit
      -- CP-element group 839: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Sample/ra
      -- 
    ra_11913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 839_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_2675_inst_ack_0, ack => minSumDecode_CP_6680_elements(839)); -- 
    -- CP-element group 840:  transition  input  no-bypass 
    -- CP-element group 840: predecessors 
    -- CP-element group 840: 	834 
    -- CP-element group 840: successors 
    -- CP-element group 840: 	103 
    -- CP-element group 840:  members (4) 
      -- CP-element group 840: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/$exit
      -- CP-element group 840: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_update_completed_
      -- CP-element group 840: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Update/$exit
      -- CP-element group 840: 	 branch_block_stmt_1353/assign_stmt_2664_to_assign_stmt_2676/SLT_i32_u1_2675_Update/ca
      -- 
    ca_11918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 840_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SLT_i32_u1_2675_inst_ack_1, ack => minSumDecode_CP_6680_elements(840)); -- 
    -- CP-element group 841:  transition  bypass 
    -- CP-element group 841: predecessors 
    -- CP-element group 841: 	103 
    -- CP-element group 841: successors 
    -- CP-element group 841:  members (1) 
      -- CP-element group 841: 	 branch_block_stmt_1353/if_stmt_2677_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(841) <= minSumDecode_CP_6680_elements(103);
    -- CP-element group 842:  transition  output  bypass 
    -- CP-element group 842: predecessors 
    -- CP-element group 842: 	103 
    -- CP-element group 842: successors 
    -- CP-element group 842: 	843 
    -- CP-element group 842:  members (3) 
      -- CP-element group 842: 	 branch_block_stmt_1353/if_stmt_2677_eval_test/$entry
      -- CP-element group 842: 	 branch_block_stmt_1353/if_stmt_2677_eval_test/$exit
      -- CP-element group 842: 	 branch_block_stmt_1353/if_stmt_2677_eval_test/branch_req
      -- 
    branch_req_11926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(842), ack => if_stmt_2677_branch_req_0); -- 
    minSumDecode_CP_6680_elements(842) <= minSumDecode_CP_6680_elements(103);
    -- CP-element group 843:  branch  place  bypass 
    -- CP-element group 843: predecessors 
    -- CP-element group 843: 	842 
    -- CP-element group 843: successors 
    -- CP-element group 843: 	844 
    -- CP-element group 843: 	846 
    -- CP-element group 843:  members (1) 
      -- CP-element group 843: 	 branch_block_stmt_1353/R_iNsTr_79_2678_place
      -- 
    minSumDecode_CP_6680_elements(843) <= minSumDecode_CP_6680_elements(842);
    -- CP-element group 844:  transition  bypass 
    -- CP-element group 844: predecessors 
    -- CP-element group 844: 	843 
    -- CP-element group 844: successors 
    -- CP-element group 844: 	845 
    -- CP-element group 844:  members (1) 
      -- CP-element group 844: 	 branch_block_stmt_1353/if_stmt_2677_if_link/$entry
      -- 
    minSumDecode_CP_6680_elements(844) <= minSumDecode_CP_6680_elements(843);
    -- CP-element group 845:  transition  input  no-bypass 
    -- CP-element group 845: predecessors 
    -- CP-element group 845: 	844 
    -- CP-element group 845: successors 
    -- CP-element group 845: 	848 
    -- CP-element group 845:  members (2) 
      -- CP-element group 845: 	 branch_block_stmt_1353/if_stmt_2677_if_link/$exit
      -- CP-element group 845: 	 branch_block_stmt_1353/if_stmt_2677_if_link/if_choice_transition
      -- 
    if_choice_transition_11931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 845_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2677_branch_ack_1, ack => minSumDecode_CP_6680_elements(845)); -- 
    -- CP-element group 846:  transition  bypass 
    -- CP-element group 846: predecessors 
    -- CP-element group 846: 	843 
    -- CP-element group 846: successors 
    -- CP-element group 846: 	847 
    -- CP-element group 846:  members (1) 
      -- CP-element group 846: 	 branch_block_stmt_1353/if_stmt_2677_else_link/$entry
      -- 
    minSumDecode_CP_6680_elements(846) <= minSumDecode_CP_6680_elements(843);
    -- CP-element group 847:  transition  input  no-bypass 
    -- CP-element group 847: predecessors 
    -- CP-element group 847: 	846 
    -- CP-element group 847: successors 
    -- CP-element group 847: 	849 
    -- CP-element group 847:  members (2) 
      -- CP-element group 847: 	 branch_block_stmt_1353/if_stmt_2677_else_link/$exit
      -- CP-element group 847: 	 branch_block_stmt_1353/if_stmt_2677_else_link/else_choice_transition
      -- 
    else_choice_transition_11935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 847_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2677_branch_ack_0, ack => minSumDecode_CP_6680_elements(847)); -- 
    -- CP-element group 848:  place  bypass 
    -- CP-element group 848: predecessors 
    -- CP-element group 848: 	845 
    -- CP-element group 848: successors 
    -- CP-element group 848: 	1202 
    -- CP-element group 848:  members (1) 
      -- CP-element group 848: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13
      -- 
    minSumDecode_CP_6680_elements(848) <= minSumDecode_CP_6680_elements(845);
    -- CP-element group 849:  place  bypass 
    -- CP-element group 849: predecessors 
    -- CP-element group 849: 	847 
    -- CP-element group 849: successors 
    -- CP-element group 849: 	1212 
    -- CP-element group 849:  members (1) 
      -- CP-element group 849: 	 branch_block_stmt_1353/bbx_xnphx_xi13_send_outputx_xexitx_xloopexit
      -- 
    minSumDecode_CP_6680_elements(849) <= minSumDecode_CP_6680_elements(847);
    -- CP-element group 850:  fork  transition  output  bypass 
    -- CP-element group 850: predecessors 
    -- CP-element group 850: 	104 
    -- CP-element group 850: successors 
    -- CP-element group 850: 	851 
    -- CP-element group 850: 	852 
    -- CP-element group 850:  members (13) 
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_root_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_update_start_
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/word_0/rr
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_word_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/word_0/cr
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/$entry
      -- CP-element group 850: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/$entry
      -- 
    cr_11967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(850), ack => LOAD_Nitr_required_2685_load_0_req_1); -- 
    rr_11956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(850), ack => LOAD_Nitr_required_2685_load_0_req_0); -- 
    minSumDecode_CP_6680_elements(850) <= minSumDecode_CP_6680_elements(104);
    -- CP-element group 851:  transition  input  no-bypass 
    -- CP-element group 851: predecessors 
    -- CP-element group 851: 	850 
    -- CP-element group 851: successors 
    -- CP-element group 851:  members (5) 
      -- CP-element group 851: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/word_0/$exit
      -- CP-element group 851: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/word_0/ra
      -- CP-element group 851: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/word_access_start/$exit
      -- CP-element group 851: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Sample/$exit
      -- CP-element group 851: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_sample_completed_
      -- 
    ra_11957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 851_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_Nitr_required_2685_load_0_ack_0, ack => minSumDecode_CP_6680_elements(851)); -- 
    -- CP-element group 852:  transition  input  no-bypass 
    -- CP-element group 852: predecessors 
    -- CP-element group 852: 	850 
    -- CP-element group 852: successors 
    -- CP-element group 852: 	105 
    -- CP-element group 852:  members (10) 
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_update_completed_
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/$exit
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/$exit
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/LOAD_Nitr_required_2685_Merge/$entry
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/word_0/ca
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/$exit
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/word_access_complete/word_0/$exit
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/LOAD_Nitr_required_2685_Merge/$exit
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/LOAD_Nitr_required_2685_Merge/merge_req
      -- CP-element group 852: 	 branch_block_stmt_1353/assign_stmt_2686/LOAD_Nitr_required_2685_Update/LOAD_Nitr_required_2685_Merge/merge_ack
      -- 
    ca_11968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 852_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_Nitr_required_2685_load_0_ack_1, ack => minSumDecode_CP_6680_elements(852)); -- 
    -- CP-element group 853:  transition  output  bypass 
    -- CP-element group 853: predecessors 
    -- CP-element group 853: 	106 
    -- CP-element group 853: successors 
    -- CP-element group 853: 	854 
    -- CP-element group 853:  members (4) 
      -- CP-element group 853: 	 branch_block_stmt_1353/assign_stmt_2700/$entry
      -- CP-element group 853: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_sample_start_
      -- CP-element group 853: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Sample/$entry
      -- CP-element group 853: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Sample/req
      -- 
    req_11984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(853), ack => WPIPE_nitr_required_2698_inst_req_0); -- 
    minSumDecode_CP_6680_elements(853) <= minSumDecode_CP_6680_elements(106);
    -- CP-element group 854:  transition  input  output  no-bypass 
    -- CP-element group 854: predecessors 
    -- CP-element group 854: 	853 
    -- CP-element group 854: successors 
    -- CP-element group 854: 	855 
    -- CP-element group 854:  members (6) 
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_sample_completed_
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_update_start_
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Sample/$exit
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Sample/ack
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Update/$entry
      -- CP-element group 854: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Update/req
      -- 
    ack_11985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 854_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nitr_required_2698_inst_ack_0, ack => minSumDecode_CP_6680_elements(854)); -- 
    req_11989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(854), ack => WPIPE_nitr_required_2698_inst_req_1); -- 
    -- CP-element group 855:  transition  input  no-bypass 
    -- CP-element group 855: predecessors 
    -- CP-element group 855: 	854 
    -- CP-element group 855: successors 
    -- CP-element group 855: 	107 
    -- CP-element group 855:  members (4) 
      -- CP-element group 855: 	 branch_block_stmt_1353/assign_stmt_2700/$exit
      -- CP-element group 855: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_update_completed_
      -- CP-element group 855: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Update/$exit
      -- CP-element group 855: 	 branch_block_stmt_1353/assign_stmt_2700/WPIPE_nitr_required_2698_Update/ack
      -- 
    ack_11990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 855_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nitr_required_2698_inst_ack_1, ack => minSumDecode_CP_6680_elements(855)); -- 
    -- CP-element group 856:  transition  bypass 
    -- CP-element group 856: predecessors 
    -- CP-element group 856: 	1 
    -- CP-element group 856: successors 
    -- CP-element group 856: 	858 
    -- CP-element group 856:  members (2) 
      -- CP-element group 856: 	 branch_block_stmt_1353/bb_0_bb_1_PhiReq/$entry
      -- CP-element group 856: 	 branch_block_stmt_1353/bb_0_bb_1_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(856) <= minSumDecode_CP_6680_elements(1);
    -- CP-element group 857:  transition  bypass 
    -- CP-element group 857: predecessors 
    -- CP-element group 857: 	107 
    -- CP-element group 857: successors 
    -- CP-element group 857: 	858 
    -- CP-element group 857:  members (2) 
      -- CP-element group 857: 	 branch_block_stmt_1353/send_outputx_xexit_bb_1_PhiReq/$entry
      -- CP-element group 857: 	 branch_block_stmt_1353/send_outputx_xexit_bb_1_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(857) <= minSumDecode_CP_6680_elements(107);
    -- CP-element group 858:  merge  place  bypass 
    -- CP-element group 858: predecessors 
    -- CP-element group 858: 	856 
    -- CP-element group 858: 	857 
    -- CP-element group 858: successors 
    -- CP-element group 858: 	859 
    -- CP-element group 858:  members (1) 
      -- CP-element group 858: 	 branch_block_stmt_1353/merge_stmt_1355_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(858) <= OrReduce(minSumDecode_CP_6680_elements(856) & minSumDecode_CP_6680_elements(857));
    -- CP-element group 859:  transition  bypass 
    -- CP-element group 859: predecessors 
    -- CP-element group 859: 	858 
    -- CP-element group 859: successors 
    -- CP-element group 859: 	3 
    -- CP-element group 859:  members (3) 
      -- CP-element group 859: 	 branch_block_stmt_1353/merge_stmt_1355_PhiAck/$entry
      -- CP-element group 859: 	 branch_block_stmt_1353/merge_stmt_1355_PhiAck/$exit
      -- CP-element group 859: 	 branch_block_stmt_1353/merge_stmt_1355_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(859) <= minSumDecode_CP_6680_elements(858);
    -- CP-element group 860:  transition  bypass 
    -- CP-element group 860: predecessors 
    -- CP-element group 860: 	124 
    -- CP-element group 860: successors 
    -- CP-element group 860: 	861 
    -- CP-element group 860:  members (2) 
      -- CP-element group 860: 	 branch_block_stmt_1353/bb_1_bbx_xnphx_xix_xpreheader_PhiReq/$entry
      -- CP-element group 860: 	 branch_block_stmt_1353/bb_1_bbx_xnphx_xix_xpreheader_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(860) <= minSumDecode_CP_6680_elements(124);
    -- CP-element group 861:  place  bypass 
    -- CP-element group 861: predecessors 
    -- CP-element group 861: 	860 
    -- CP-element group 861: successors 
    -- CP-element group 861: 	862 
    -- CP-element group 861:  members (1) 
      -- CP-element group 861: 	 branch_block_stmt_1353/merge_stmt_1372_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(861) <= minSumDecode_CP_6680_elements(860);
    -- CP-element group 862:  transition  bypass 
    -- CP-element group 862: predecessors 
    -- CP-element group 862: 	861 
    -- CP-element group 862: successors 
    -- CP-element group 862: 	6 
    -- CP-element group 862:  members (3) 
      -- CP-element group 862: 	 branch_block_stmt_1353/merge_stmt_1372_PhiAck/$entry
      -- CP-element group 862: 	 branch_block_stmt_1353/merge_stmt_1372_PhiAck/$exit
      -- CP-element group 862: 	 branch_block_stmt_1353/merge_stmt_1372_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(862) <= minSumDecode_CP_6680_elements(861);
    -- CP-element group 863:  transition  bypass 
    -- CP-element group 863: predecessors 
    -- CP-element group 863: 	6 
    -- CP-element group 863: successors 
    -- CP-element group 863: 	864 
    -- CP-element group 863:  members (3) 
      -- CP-element group 863: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 863: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/$entry
      -- CP-element group 863: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(863) <= minSumDecode_CP_6680_elements(6);
    -- CP-element group 864:  transition  bypass 
    -- CP-element group 864: predecessors 
    -- CP-element group 864: 	863 
    -- CP-element group 864: successors 
    -- CP-element group 864: 	865 
    -- CP-element group 864:  members (1) 
      -- CP-element group 864: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1379_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(864) is a control-delay.
    cp_element_864_delay: control_delay_element  generic map(name => " 864_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(863), ack => minSumDecode_CP_6680_elements(864), clk => clk, reset =>reset);
    -- CP-element group 865:  transition  output  bypass 
    -- CP-element group 865: predecessors 
    -- CP-element group 865: 	864 
    -- CP-element group 865: successors 
    -- CP-element group 865: 	866 
    -- CP-element group 865:  members (4) 
      -- CP-element group 865: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 865: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/$exit
      -- CP-element group 865: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$exit
      -- CP-element group 865: 	 branch_block_stmt_1353/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_1375/phi_stmt_1375_req
      -- 
    phi_stmt_1375_req_12024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1375_req_12024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(865), ack => phi_stmt_1375_req_0); -- 
    minSumDecode_CP_6680_elements(865) <= minSumDecode_CP_6680_elements(864);
    -- CP-element group 866:  place  bypass 
    -- CP-element group 866: predecessors 
    -- CP-element group 866: 	865 
    -- CP-element group 866: successors 
    -- CP-element group 866: 	867 
    -- CP-element group 866:  members (1) 
      -- CP-element group 866: 	 branch_block_stmt_1353/merge_stmt_1374_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(866) <= minSumDecode_CP_6680_elements(865);
    -- CP-element group 867:  transition  bypass 
    -- CP-element group 867: predecessors 
    -- CP-element group 867: 	866 
    -- CP-element group 867: successors 
    -- CP-element group 867: 	868 
    -- CP-element group 867:  members (1) 
      -- CP-element group 867: 	 branch_block_stmt_1353/merge_stmt_1374_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(867) <= minSumDecode_CP_6680_elements(866);
    -- CP-element group 868:  transition  input  no-bypass 
    -- CP-element group 868: predecessors 
    -- CP-element group 868: 	867 
    -- CP-element group 868: successors 
    -- CP-element group 868: 	7 
    -- CP-element group 868:  members (2) 
      -- CP-element group 868: 	 branch_block_stmt_1353/merge_stmt_1374_PhiAck/$exit
      -- CP-element group 868: 	 branch_block_stmt_1353/merge_stmt_1374_PhiAck/phi_stmt_1375_ack
      -- 
    phi_stmt_1375_ack_12029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 868_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1375_ack_0, ack => minSumDecode_CP_6680_elements(868)); -- 
    -- CP-element group 869:  transition  bypass 
    -- CP-element group 869: predecessors 
    -- CP-element group 869: 	9 
    -- CP-element group 869: successors 
    -- CP-element group 869:  members (1) 
      -- CP-element group 869: 	 branch_block_stmt_1353/merge_stmt_1443_dead_link/$entry
      -- 
    minSumDecode_CP_6680_elements(869) <= minSumDecode_CP_6680_elements(9);
    -- CP-element group 870:  fork  transition  output  bypass 
    -- CP-element group 870: predecessors 
    -- CP-element group 870: 	214 
    -- CP-element group 870: successors 
    -- CP-element group 870: 	871 
    -- CP-element group 870: 	872 
    -- CP-element group 870:  members (9) 
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Sample/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Sample/rr
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Update/$entry
      -- CP-element group 870: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Update/cr
      -- 
    rr_12052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(870), ack => type_cast_1447_inst_req_0); -- 
    cr_12057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(870), ack => type_cast_1447_inst_req_1); -- 
    minSumDecode_CP_6680_elements(870) <= minSumDecode_CP_6680_elements(214);
    -- CP-element group 871:  transition  input  no-bypass 
    -- CP-element group 871: predecessors 
    -- CP-element group 871: 	870 
    -- CP-element group 871: successors 
    -- CP-element group 871: 	873 
    -- CP-element group 871:  members (2) 
      -- CP-element group 871: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Sample/$exit
      -- CP-element group 871: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Sample/ra
      -- 
    ra_12053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 871_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_0, ack => minSumDecode_CP_6680_elements(871)); -- 
    -- CP-element group 872:  transition  input  no-bypass 
    -- CP-element group 872: predecessors 
    -- CP-element group 872: 	870 
    -- CP-element group 872: successors 
    -- CP-element group 872: 	873 
    -- CP-element group 872:  members (2) 
      -- CP-element group 872: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Update/$exit
      -- CP-element group 872: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/Update/ca
      -- 
    ca_12058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 872_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_1, ack => minSumDecode_CP_6680_elements(872)); -- 
    -- CP-element group 873:  join  transition  output  bypass 
    -- CP-element group 873: predecessors 
    -- CP-element group 873: 	871 
    -- CP-element group 873: 	872 
    -- CP-element group 873: successors 
    -- CP-element group 873: 	874 
    -- CP-element group 873:  members (6) 
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/$exit
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/$exit
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/$exit
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/$exit
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_sources/type_cast_1447/SplitProtocol/$exit
      -- CP-element group 873: 	 branch_block_stmt_1353/bbx_xnphx_xi_readCodeBlockx_xexit_PhiReq/phi_stmt_1444/phi_stmt_1444_req
      -- 
    phi_stmt_1444_req_12059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1444_req_12059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(873), ack => phi_stmt_1444_req_0); -- 
    minSumDecode_cp_element_group_873: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_873"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(871) & minSumDecode_CP_6680_elements(872);
      gj_minSumDecode_cp_element_group_873 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(873), clk => clk, reset => reset); --
    end block;
    -- CP-element group 874:  place  bypass 
    -- CP-element group 874: predecessors 
    -- CP-element group 874: 	873 
    -- CP-element group 874: successors 
    -- CP-element group 874: 	875 
    -- CP-element group 874:  members (1) 
      -- CP-element group 874: 	 branch_block_stmt_1353/merge_stmt_1443_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(874) <= minSumDecode_CP_6680_elements(873);
    -- CP-element group 875:  transition  bypass 
    -- CP-element group 875: predecessors 
    -- CP-element group 875: 	874 
    -- CP-element group 875: successors 
    -- CP-element group 875: 	876 
    -- CP-element group 875:  members (1) 
      -- CP-element group 875: 	 branch_block_stmt_1353/merge_stmt_1443_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(875) <= minSumDecode_CP_6680_elements(874);
    -- CP-element group 876:  transition  input  no-bypass 
    -- CP-element group 876: predecessors 
    -- CP-element group 876: 	875 
    -- CP-element group 876: successors 
    -- CP-element group 876: 	10 
    -- CP-element group 876:  members (2) 
      -- CP-element group 876: 	 branch_block_stmt_1353/merge_stmt_1443_PhiAck/$exit
      -- CP-element group 876: 	 branch_block_stmt_1353/merge_stmt_1443_PhiAck/phi_stmt_1444_ack
      -- 
    phi_stmt_1444_ack_12064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 876_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1444_ack_0, ack => minSumDecode_CP_6680_elements(876)); -- 
    -- CP-element group 877:  transition  bypass 
    -- CP-element group 877: predecessors 
    -- CP-element group 877: 	226 
    -- CP-element group 877: successors 
    -- CP-element group 877: 	878 
    -- CP-element group 877:  members (2) 
      -- CP-element group 877: 	 branch_block_stmt_1353/readCodeBlockx_xexit_bbx_xnphx_xi1_PhiReq/$entry
      -- CP-element group 877: 	 branch_block_stmt_1353/readCodeBlockx_xexit_bbx_xnphx_xi1_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(877) <= minSumDecode_CP_6680_elements(226);
    -- CP-element group 878:  place  bypass 
    -- CP-element group 878: predecessors 
    -- CP-element group 878: 	877 
    -- CP-element group 878: successors 
    -- CP-element group 878: 	879 
    -- CP-element group 878:  members (1) 
      -- CP-element group 878: 	 branch_block_stmt_1353/merge_stmt_1461_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(878) <= minSumDecode_CP_6680_elements(877);
    -- CP-element group 879:  transition  bypass 
    -- CP-element group 879: predecessors 
    -- CP-element group 879: 	878 
    -- CP-element group 879: successors 
    -- CP-element group 879: 	12 
    -- CP-element group 879:  members (3) 
      -- CP-element group 879: 	 branch_block_stmt_1353/merge_stmt_1461_PhiAck/$entry
      -- CP-element group 879: 	 branch_block_stmt_1353/merge_stmt_1461_PhiAck/$exit
      -- CP-element group 879: 	 branch_block_stmt_1353/merge_stmt_1461_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(879) <= minSumDecode_CP_6680_elements(878);
    -- CP-element group 880:  fork  transition  output  bypass 
    -- CP-element group 880: predecessors 
    -- CP-element group 880: 	274 
    -- CP-element group 880: successors 
    -- CP-element group 880: 	881 
    -- CP-element group 880: 	882 
    -- CP-element group 880:  members (9) 
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/rr
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/$entry
      -- CP-element group 880: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/cr
      -- 
    rr_12095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(880), ack => type_cast_1510_inst_req_0); -- 
    cr_12100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(880), ack => type_cast_1510_inst_req_1); -- 
    minSumDecode_CP_6680_elements(880) <= minSumDecode_CP_6680_elements(274);
    -- CP-element group 881:  transition  input  no-bypass 
    -- CP-element group 881: predecessors 
    -- CP-element group 881: 	880 
    -- CP-element group 881: successors 
    -- CP-element group 881: 	883 
    -- CP-element group 881:  members (2) 
      -- CP-element group 881: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/$exit
      -- CP-element group 881: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Sample/ra
      -- 
    ra_12096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 881_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_0, ack => minSumDecode_CP_6680_elements(881)); -- 
    -- CP-element group 882:  transition  input  no-bypass 
    -- CP-element group 882: predecessors 
    -- CP-element group 882: 	880 
    -- CP-element group 882: successors 
    -- CP-element group 882: 	883 
    -- CP-element group 882:  members (2) 
      -- CP-element group 882: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/$exit
      -- CP-element group 882: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/Update/ca
      -- 
    ca_12101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 882_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_1, ack => minSumDecode_CP_6680_elements(882)); -- 
    -- CP-element group 883:  join  transition  output  bypass 
    -- CP-element group 883: predecessors 
    -- CP-element group 883: 	881 
    -- CP-element group 883: 	882 
    -- CP-element group 883: successors 
    -- CP-element group 883: 	887 
    -- CP-element group 883:  members (6) 
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/$exit
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/$exit
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$exit
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/$exit
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1510/SplitProtocol/$exit
      -- CP-element group 883: 	 branch_block_stmt_1353/bb_6_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_req
      -- 
    phi_stmt_1504_req_12102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1504_req_12102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(883), ack => phi_stmt_1504_req_1); -- 
    minSumDecode_cp_element_group_883: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_883"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(881) & minSumDecode_CP_6680_elements(882);
      gj_minSumDecode_cp_element_group_883 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(883), clk => clk, reset => reset); --
    end block;
    -- CP-element group 884:  transition  bypass 
    -- CP-element group 884: predecessors 
    -- CP-element group 884: 	13 
    -- CP-element group 884: successors 
    -- CP-element group 884: 	885 
    -- CP-element group 884:  members (3) 
      -- CP-element group 884: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/$entry
      -- CP-element group 884: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/$entry
      -- CP-element group 884: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(884) <= minSumDecode_CP_6680_elements(13);
    -- CP-element group 885:  transition  bypass 
    -- CP-element group 885: predecessors 
    -- CP-element group 885: 	884 
    -- CP-element group 885: successors 
    -- CP-element group 885: 	886 
    -- CP-element group 885:  members (1) 
      -- CP-element group 885: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/type_cast_1508_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(885) is a control-delay.
    cp_element_885_delay: control_delay_element  generic map(name => " 885_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(884), ack => minSumDecode_CP_6680_elements(885), clk => clk, reset =>reset);
    -- CP-element group 886:  transition  output  bypass 
    -- CP-element group 886: predecessors 
    -- CP-element group 886: 	885 
    -- CP-element group 886: successors 
    -- CP-element group 886: 	887 
    -- CP-element group 886:  members (4) 
      -- CP-element group 886: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/$exit
      -- CP-element group 886: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/$exit
      -- CP-element group 886: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_sources/$exit
      -- CP-element group 886: 	 branch_block_stmt_1353/bbx_xnphx_xi1_bb_6_PhiReq/phi_stmt_1504/phi_stmt_1504_req
      -- 
    phi_stmt_1504_req_12113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1504_req_12113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(886), ack => phi_stmt_1504_req_0); -- 
    minSumDecode_CP_6680_elements(886) <= minSumDecode_CP_6680_elements(885);
    -- CP-element group 887:  merge  place  bypass 
    -- CP-element group 887: predecessors 
    -- CP-element group 887: 	883 
    -- CP-element group 887: 	886 
    -- CP-element group 887: successors 
    -- CP-element group 887: 	888 
    -- CP-element group 887:  members (1) 
      -- CP-element group 887: 	 branch_block_stmt_1353/merge_stmt_1503_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(887) <= OrReduce(minSumDecode_CP_6680_elements(883) & minSumDecode_CP_6680_elements(886));
    -- CP-element group 888:  transition  bypass 
    -- CP-element group 888: predecessors 
    -- CP-element group 888: 	887 
    -- CP-element group 888: successors 
    -- CP-element group 888: 	889 
    -- CP-element group 888:  members (1) 
      -- CP-element group 888: 	 branch_block_stmt_1353/merge_stmt_1503_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(888) <= minSumDecode_CP_6680_elements(887);
    -- CP-element group 889:  transition  input  no-bypass 
    -- CP-element group 889: predecessors 
    -- CP-element group 889: 	888 
    -- CP-element group 889: successors 
    -- CP-element group 889: 	14 
    -- CP-element group 889:  members (2) 
      -- CP-element group 889: 	 branch_block_stmt_1353/merge_stmt_1503_PhiAck/$exit
      -- CP-element group 889: 	 branch_block_stmt_1353/merge_stmt_1503_PhiAck/phi_stmt_1504_ack
      -- 
    phi_stmt_1504_ack_12118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 889_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1504_ack_0, ack => minSumDecode_CP_6680_elements(889)); -- 
    -- CP-element group 890:  transition  bypass 
    -- CP-element group 890: predecessors 
    -- CP-element group 890: 	273 
    -- CP-element group 890: successors 
    -- CP-element group 890: 	891 
    -- CP-element group 890:  members (2) 
      -- CP-element group 890: 	 branch_block_stmt_1353/bb_6_initialize_aPriorix_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 890: 	 branch_block_stmt_1353/bb_6_initialize_aPriorix_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(890) <= minSumDecode_CP_6680_elements(273);
    -- CP-element group 891:  place  bypass 
    -- CP-element group 891: predecessors 
    -- CP-element group 891: 	890 
    -- CP-element group 891: successors 
    -- CP-element group 891: 	892 
    -- CP-element group 891:  members (1) 
      -- CP-element group 891: 	 branch_block_stmt_1353/merge_stmt_1558_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(891) <= minSumDecode_CP_6680_elements(890);
    -- CP-element group 892:  transition  bypass 
    -- CP-element group 892: predecessors 
    -- CP-element group 892: 	891 
    -- CP-element group 892: successors 
    -- CP-element group 892: 	16 
    -- CP-element group 892:  members (3) 
      -- CP-element group 892: 	 branch_block_stmt_1353/merge_stmt_1558_PhiAck/$entry
      -- CP-element group 892: 	 branch_block_stmt_1353/merge_stmt_1558_PhiAck/$exit
      -- CP-element group 892: 	 branch_block_stmt_1353/merge_stmt_1558_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(892) <= minSumDecode_CP_6680_elements(891);
    -- CP-element group 893:  transition  bypass 
    -- CP-element group 893: predecessors 
    -- CP-element group 893: 	123 
    -- CP-element group 893: successors 
    -- CP-element group 893: 	894 
    -- CP-element group 893:  members (3) 
      -- CP-element group 893: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/$entry
      -- CP-element group 893: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$entry
      -- CP-element group 893: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(893) <= minSumDecode_CP_6680_elements(123);
    -- CP-element group 894:  transition  bypass 
    -- CP-element group 894: predecessors 
    -- CP-element group 894: 	893 
    -- CP-element group 894: successors 
    -- CP-element group 894: 	895 
    -- CP-element group 894:  members (1) 
      -- CP-element group 894: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1565_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(894) is a control-delay.
    cp_element_894_delay: control_delay_element  generic map(name => " 894_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(893), ack => minSumDecode_CP_6680_elements(894), clk => clk, reset =>reset);
    -- CP-element group 895:  transition  output  bypass 
    -- CP-element group 895: predecessors 
    -- CP-element group 895: 	894 
    -- CP-element group 895: successors 
    -- CP-element group 895: 	903 
    -- CP-element group 895:  members (4) 
      -- CP-element group 895: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/$exit
      -- CP-element group 895: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$exit
      -- CP-element group 895: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$exit
      -- CP-element group 895: 	 branch_block_stmt_1353/bb_1_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_req
      -- 
    phi_stmt_1561_req_12141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1561_req_12141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(895), ack => phi_stmt_1561_req_0); -- 
    minSumDecode_CP_6680_elements(895) <= minSumDecode_CP_6680_elements(894);
    -- CP-element group 896:  fork  transition  output  bypass 
    -- CP-element group 896: predecessors 
    -- CP-element group 896: 	16 
    -- CP-element group 896: successors 
    -- CP-element group 896: 	897 
    -- CP-element group 896: 	898 
    -- CP-element group 896:  members (9) 
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Sample/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Sample/rr
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Update/$entry
      -- CP-element group 896: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Update/cr
      -- 
    rr_12160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(896), ack => type_cast_1570_inst_req_0); -- 
    cr_12165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(896), ack => type_cast_1570_inst_req_1); -- 
    minSumDecode_CP_6680_elements(896) <= minSumDecode_CP_6680_elements(16);
    -- CP-element group 897:  transition  input  no-bypass 
    -- CP-element group 897: predecessors 
    -- CP-element group 897: 	896 
    -- CP-element group 897: successors 
    -- CP-element group 897: 	899 
    -- CP-element group 897:  members (2) 
      -- CP-element group 897: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Sample/$exit
      -- CP-element group 897: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Sample/ra
      -- 
    ra_12161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 897_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_0, ack => minSumDecode_CP_6680_elements(897)); -- 
    -- CP-element group 898:  transition  input  no-bypass 
    -- CP-element group 898: predecessors 
    -- CP-element group 898: 	896 
    -- CP-element group 898: successors 
    -- CP-element group 898: 	899 
    -- CP-element group 898:  members (2) 
      -- CP-element group 898: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Update/$exit
      -- CP-element group 898: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/Update/ca
      -- 
    ca_12166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 898_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_1, ack => minSumDecode_CP_6680_elements(898)); -- 
    -- CP-element group 899:  join  transition  output  bypass 
    -- CP-element group 899: predecessors 
    -- CP-element group 899: 	897 
    -- CP-element group 899: 	898 
    -- CP-element group 899: successors 
    -- CP-element group 899: 	903 
    -- CP-element group 899:  members (6) 
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/$exit
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$exit
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$exit
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/$exit
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1570/SplitProtocol/$exit
      -- CP-element group 899: 	 branch_block_stmt_1353/initialize_aPriorix_xexitx_xloopexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_req
      -- 
    phi_stmt_1561_req_12167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1561_req_12167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(899), ack => phi_stmt_1561_req_2); -- 
    minSumDecode_cp_element_group_899: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_899"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(897) & minSumDecode_CP_6680_elements(898);
      gj_minSumDecode_cp_element_group_899 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(899), clk => clk, reset => reset); --
    end block;
    -- CP-element group 900:  transition  bypass 
    -- CP-element group 900: predecessors 
    -- CP-element group 900: 	225 
    -- CP-element group 900: successors 
    -- CP-element group 900: 	901 
    -- CP-element group 900:  members (3) 
      -- CP-element group 900: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/$entry
      -- CP-element group 900: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$entry
      -- CP-element group 900: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(900) <= minSumDecode_CP_6680_elements(225);
    -- CP-element group 901:  transition  bypass 
    -- CP-element group 901: predecessors 
    -- CP-element group 901: 	900 
    -- CP-element group 901: successors 
    -- CP-element group 901: 	902 
    -- CP-element group 901:  members (1) 
      -- CP-element group 901: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1568_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(901) is a control-delay.
    cp_element_901_delay: control_delay_element  generic map(name => " 901_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(900), ack => minSumDecode_CP_6680_elements(901), clk => clk, reset =>reset);
    -- CP-element group 902:  transition  output  bypass 
    -- CP-element group 902: predecessors 
    -- CP-element group 902: 	901 
    -- CP-element group 902: successors 
    -- CP-element group 902: 	903 
    -- CP-element group 902:  members (4) 
      -- CP-element group 902: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/$exit
      -- CP-element group 902: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/$exit
      -- CP-element group 902: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$exit
      -- CP-element group 902: 	 branch_block_stmt_1353/readCodeBlockx_xexit_initialize_aPriorix_xexit_PhiReq/phi_stmt_1561/phi_stmt_1561_req
      -- 
    phi_stmt_1561_req_12178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1561_req_12178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(902), ack => phi_stmt_1561_req_1); -- 
    minSumDecode_CP_6680_elements(902) <= minSumDecode_CP_6680_elements(901);
    -- CP-element group 903:  merge  place  bypass 
    -- CP-element group 903: predecessors 
    -- CP-element group 903: 	895 
    -- CP-element group 903: 	899 
    -- CP-element group 903: 	902 
    -- CP-element group 903: successors 
    -- CP-element group 903: 	904 
    -- CP-element group 903:  members (1) 
      -- CP-element group 903: 	 branch_block_stmt_1353/merge_stmt_1560_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(903) <= OrReduce(minSumDecode_CP_6680_elements(895) & minSumDecode_CP_6680_elements(899) & minSumDecode_CP_6680_elements(902));
    -- CP-element group 904:  transition  bypass 
    -- CP-element group 904: predecessors 
    -- CP-element group 904: 	903 
    -- CP-element group 904: successors 
    -- CP-element group 904: 	905 
    -- CP-element group 904:  members (1) 
      -- CP-element group 904: 	 branch_block_stmt_1353/merge_stmt_1560_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(904) <= minSumDecode_CP_6680_elements(903);
    -- CP-element group 905:  transition  input  no-bypass 
    -- CP-element group 905: predecessors 
    -- CP-element group 905: 	904 
    -- CP-element group 905: successors 
    -- CP-element group 905: 	17 
    -- CP-element group 905:  members (2) 
      -- CP-element group 905: 	 branch_block_stmt_1353/merge_stmt_1560_PhiAck/$exit
      -- CP-element group 905: 	 branch_block_stmt_1353/merge_stmt_1560_PhiAck/phi_stmt_1561_ack
      -- 
    phi_stmt_1561_ack_12183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 905_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1561_ack_0, ack => minSumDecode_CP_6680_elements(905)); -- 
    -- CP-element group 906:  transition  bypass 
    -- CP-element group 906: predecessors 
    -- CP-element group 906: 	288 
    -- CP-element group 906: successors 
    -- CP-element group 906: 	907 
    -- CP-element group 906:  members (2) 
      -- CP-element group 906: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_bbx_xnphx_xi5_PhiReq/$entry
      -- CP-element group 906: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_bbx_xnphx_xi5_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(906) <= minSumDecode_CP_6680_elements(288);
    -- CP-element group 907:  place  bypass 
    -- CP-element group 907: predecessors 
    -- CP-element group 907: 	906 
    -- CP-element group 907: successors 
    -- CP-element group 907: 	908 
    -- CP-element group 907:  members (1) 
      -- CP-element group 907: 	 branch_block_stmt_1353/merge_stmt_1587_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(907) <= minSumDecode_CP_6680_elements(906);
    -- CP-element group 908:  transition  bypass 
    -- CP-element group 908: predecessors 
    -- CP-element group 908: 	907 
    -- CP-element group 908: successors 
    -- CP-element group 908: 	19 
    -- CP-element group 908:  members (3) 
      -- CP-element group 908: 	 branch_block_stmt_1353/merge_stmt_1587_PhiAck/$entry
      -- CP-element group 908: 	 branch_block_stmt_1353/merge_stmt_1587_PhiAck/$exit
      -- CP-element group 908: 	 branch_block_stmt_1353/merge_stmt_1587_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(908) <= minSumDecode_CP_6680_elements(907);
    -- CP-element group 909:  fork  transition  output  bypass 
    -- CP-element group 909: predecessors 
    -- CP-element group 909: 	335 
    -- CP-element group 909: successors 
    -- CP-element group 909: 	910 
    -- CP-element group 909: 	911 
    -- CP-element group 909:  members (9) 
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/rr
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/$entry
      -- CP-element group 909: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/cr
      -- 
    rr_12214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(909), ack => type_cast_1625_inst_req_0); -- 
    cr_12219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(909), ack => type_cast_1625_inst_req_1); -- 
    minSumDecode_CP_6680_elements(909) <= minSumDecode_CP_6680_elements(335);
    -- CP-element group 910:  transition  input  no-bypass 
    -- CP-element group 910: predecessors 
    -- CP-element group 910: 	909 
    -- CP-element group 910: successors 
    -- CP-element group 910: 	912 
    -- CP-element group 910:  members (2) 
      -- CP-element group 910: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/$exit
      -- CP-element group 910: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Sample/ra
      -- 
    ra_12215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 910_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => minSumDecode_CP_6680_elements(910)); -- 
    -- CP-element group 911:  transition  input  no-bypass 
    -- CP-element group 911: predecessors 
    -- CP-element group 911: 	909 
    -- CP-element group 911: successors 
    -- CP-element group 911: 	912 
    -- CP-element group 911:  members (2) 
      -- CP-element group 911: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/$exit
      -- CP-element group 911: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/Update/ca
      -- 
    ca_12220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 911_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => minSumDecode_CP_6680_elements(911)); -- 
    -- CP-element group 912:  join  transition  output  bypass 
    -- CP-element group 912: predecessors 
    -- CP-element group 912: 	910 
    -- CP-element group 912: 	911 
    -- CP-element group 912: successors 
    -- CP-element group 912: 	916 
    -- CP-element group 912:  members (6) 
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/$exit
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/$exit
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$exit
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/$exit
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1625/SplitProtocol/$exit
      -- CP-element group 912: 	 branch_block_stmt_1353/bb_10_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_req
      -- 
    phi_stmt_1619_req_12221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1619_req_12221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(912), ack => phi_stmt_1619_req_1); -- 
    minSumDecode_cp_element_group_912: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_912"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(910) & minSumDecode_CP_6680_elements(911);
      gj_minSumDecode_cp_element_group_912 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(912), clk => clk, reset => reset); --
    end block;
    -- CP-element group 913:  transition  bypass 
    -- CP-element group 913: predecessors 
    -- CP-element group 913: 	20 
    -- CP-element group 913: successors 
    -- CP-element group 913: 	914 
    -- CP-element group 913:  members (3) 
      -- CP-element group 913: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/$entry
      -- CP-element group 913: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/$entry
      -- CP-element group 913: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(913) <= minSumDecode_CP_6680_elements(20);
    -- CP-element group 914:  transition  bypass 
    -- CP-element group 914: predecessors 
    -- CP-element group 914: 	913 
    -- CP-element group 914: successors 
    -- CP-element group 914: 	915 
    -- CP-element group 914:  members (1) 
      -- CP-element group 914: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/type_cast_1623_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(914) is a control-delay.
    cp_element_914_delay: control_delay_element  generic map(name => " 914_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(913), ack => minSumDecode_CP_6680_elements(914), clk => clk, reset =>reset);
    -- CP-element group 915:  transition  output  bypass 
    -- CP-element group 915: predecessors 
    -- CP-element group 915: 	914 
    -- CP-element group 915: successors 
    -- CP-element group 915: 	916 
    -- CP-element group 915:  members (4) 
      -- CP-element group 915: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/$exit
      -- CP-element group 915: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/$exit
      -- CP-element group 915: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_sources/$exit
      -- CP-element group 915: 	 branch_block_stmt_1353/bbx_xnphx_xi5_bb_10_PhiReq/phi_stmt_1619/phi_stmt_1619_req
      -- 
    phi_stmt_1619_req_12232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1619_req_12232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(915), ack => phi_stmt_1619_req_0); -- 
    minSumDecode_CP_6680_elements(915) <= minSumDecode_CP_6680_elements(914);
    -- CP-element group 916:  merge  place  bypass 
    -- CP-element group 916: predecessors 
    -- CP-element group 916: 	912 
    -- CP-element group 916: 	915 
    -- CP-element group 916: successors 
    -- CP-element group 916: 	917 
    -- CP-element group 916:  members (1) 
      -- CP-element group 916: 	 branch_block_stmt_1353/merge_stmt_1618_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(916) <= OrReduce(minSumDecode_CP_6680_elements(912) & minSumDecode_CP_6680_elements(915));
    -- CP-element group 917:  transition  bypass 
    -- CP-element group 917: predecessors 
    -- CP-element group 917: 	916 
    -- CP-element group 917: successors 
    -- CP-element group 917: 	918 
    -- CP-element group 917:  members (1) 
      -- CP-element group 917: 	 branch_block_stmt_1353/merge_stmt_1618_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(917) <= minSumDecode_CP_6680_elements(916);
    -- CP-element group 918:  transition  input  no-bypass 
    -- CP-element group 918: predecessors 
    -- CP-element group 918: 	917 
    -- CP-element group 918: successors 
    -- CP-element group 918: 	21 
    -- CP-element group 918:  members (2) 
      -- CP-element group 918: 	 branch_block_stmt_1353/merge_stmt_1618_PhiAck/$exit
      -- CP-element group 918: 	 branch_block_stmt_1353/merge_stmt_1618_PhiAck/phi_stmt_1619_ack
      -- 
    phi_stmt_1619_ack_12237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 918_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1619_ack_0, ack => minSumDecode_CP_6680_elements(918)); -- 
    -- CP-element group 919:  transition  bypass 
    -- CP-element group 919: predecessors 
    -- CP-element group 919: 	334 
    -- CP-element group 919: successors 
    -- CP-element group 919: 	920 
    -- CP-element group 919:  members (2) 
      -- CP-element group 919: 	 branch_block_stmt_1353/bb_10_initializeMessagex_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 919: 	 branch_block_stmt_1353/bb_10_initializeMessagex_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(919) <= minSumDecode_CP_6680_elements(334);
    -- CP-element group 920:  place  bypass 
    -- CP-element group 920: predecessors 
    -- CP-element group 920: 	919 
    -- CP-element group 920: successors 
    -- CP-element group 920: 	921 
    -- CP-element group 920:  members (1) 
      -- CP-element group 920: 	 branch_block_stmt_1353/merge_stmt_1687_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(920) <= minSumDecode_CP_6680_elements(919);
    -- CP-element group 921:  transition  bypass 
    -- CP-element group 921: predecessors 
    -- CP-element group 921: 	920 
    -- CP-element group 921: successors 
    -- CP-element group 921: 	23 
    -- CP-element group 921:  members (3) 
      -- CP-element group 921: 	 branch_block_stmt_1353/merge_stmt_1687_PhiAck/$entry
      -- CP-element group 921: 	 branch_block_stmt_1353/merge_stmt_1687_PhiAck/$exit
      -- CP-element group 921: 	 branch_block_stmt_1353/merge_stmt_1687_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(921) <= minSumDecode_CP_6680_elements(920);
    -- CP-element group 922:  fork  transition  output  bypass 
    -- CP-element group 922: predecessors 
    -- CP-element group 922: 	23 
    -- CP-element group 922: successors 
    -- CP-element group 922: 	923 
    -- CP-element group 922: 	924 
    -- CP-element group 922:  members (9) 
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Sample/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Sample/rr
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Update/$entry
      -- CP-element group 922: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Update/cr
      -- 
    rr_12268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(922), ack => type_cast_1693_inst_req_0); -- 
    cr_12273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(922), ack => type_cast_1693_inst_req_1); -- 
    minSumDecode_CP_6680_elements(922) <= minSumDecode_CP_6680_elements(23);
    -- CP-element group 923:  transition  input  no-bypass 
    -- CP-element group 923: predecessors 
    -- CP-element group 923: 	922 
    -- CP-element group 923: successors 
    -- CP-element group 923: 	925 
    -- CP-element group 923:  members (2) 
      -- CP-element group 923: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Sample/$exit
      -- CP-element group 923: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Sample/ra
      -- 
    ra_12269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 923_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1693_inst_ack_0, ack => minSumDecode_CP_6680_elements(923)); -- 
    -- CP-element group 924:  transition  input  no-bypass 
    -- CP-element group 924: predecessors 
    -- CP-element group 924: 	922 
    -- CP-element group 924: successors 
    -- CP-element group 924: 	925 
    -- CP-element group 924:  members (2) 
      -- CP-element group 924: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Update/$exit
      -- CP-element group 924: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/Update/ca
      -- 
    ca_12274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 924_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1693_inst_ack_1, ack => minSumDecode_CP_6680_elements(924)); -- 
    -- CP-element group 925:  join  transition  output  bypass 
    -- CP-element group 925: predecessors 
    -- CP-element group 925: 	923 
    -- CP-element group 925: 	924 
    -- CP-element group 925: successors 
    -- CP-element group 925: 	929 
    -- CP-element group 925:  members (6) 
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/$exit
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/$exit
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$exit
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/$exit
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1693/SplitProtocol/$exit
      -- CP-element group 925: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xloopexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_req
      -- 
    phi_stmt_1690_req_12275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1690_req_12275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(925), ack => phi_stmt_1690_req_0); -- 
    minSumDecode_cp_element_group_925: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_925"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(923) & minSumDecode_CP_6680_elements(924);
      gj_minSumDecode_cp_element_group_925 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 926:  transition  bypass 
    -- CP-element group 926: predecessors 
    -- CP-element group 926: 	287 
    -- CP-element group 926: successors 
    -- CP-element group 926: 	927 
    -- CP-element group 926:  members (3) 
      -- CP-element group 926: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/$entry
      -- CP-element group 926: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/$entry
      -- CP-element group 926: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(926) <= minSumDecode_CP_6680_elements(287);
    -- CP-element group 927:  transition  bypass 
    -- CP-element group 927: predecessors 
    -- CP-element group 927: 	926 
    -- CP-element group 927: successors 
    -- CP-element group 927: 	928 
    -- CP-element group 927:  members (1) 
      -- CP-element group 927: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/type_cast_1696_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(927) is a control-delay.
    cp_element_927_delay: control_delay_element  generic map(name => " 927_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(926), ack => minSumDecode_CP_6680_elements(927), clk => clk, reset =>reset);
    -- CP-element group 928:  transition  output  bypass 
    -- CP-element group 928: predecessors 
    -- CP-element group 928: 	927 
    -- CP-element group 928: successors 
    -- CP-element group 928: 	929 
    -- CP-element group 928:  members (4) 
      -- CP-element group 928: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/$exit
      -- CP-element group 928: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/$exit
      -- CP-element group 928: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_sources/$exit
      -- CP-element group 928: 	 branch_block_stmt_1353/initialize_aPriorix_xexit_initializeMessagex_xexitx_xpreheader_PhiReq/phi_stmt_1690/phi_stmt_1690_req
      -- 
    phi_stmt_1690_req_12286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1690_req_12286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(928), ack => phi_stmt_1690_req_1); -- 
    minSumDecode_CP_6680_elements(928) <= minSumDecode_CP_6680_elements(927);
    -- CP-element group 929:  merge  place  bypass 
    -- CP-element group 929: predecessors 
    -- CP-element group 929: 	925 
    -- CP-element group 929: 	928 
    -- CP-element group 929: successors 
    -- CP-element group 929: 	930 
    -- CP-element group 929:  members (1) 
      -- CP-element group 929: 	 branch_block_stmt_1353/merge_stmt_1689_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(929) <= OrReduce(minSumDecode_CP_6680_elements(925) & minSumDecode_CP_6680_elements(928));
    -- CP-element group 930:  transition  bypass 
    -- CP-element group 930: predecessors 
    -- CP-element group 930: 	929 
    -- CP-element group 930: successors 
    -- CP-element group 930: 	931 
    -- CP-element group 930:  members (1) 
      -- CP-element group 930: 	 branch_block_stmt_1353/merge_stmt_1689_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(930) <= minSumDecode_CP_6680_elements(929);
    -- CP-element group 931:  transition  input  no-bypass 
    -- CP-element group 931: predecessors 
    -- CP-element group 931: 	930 
    -- CP-element group 931: successors 
    -- CP-element group 931: 	24 
    -- CP-element group 931:  members (2) 
      -- CP-element group 931: 	 branch_block_stmt_1353/merge_stmt_1689_PhiAck/$exit
      -- CP-element group 931: 	 branch_block_stmt_1353/merge_stmt_1689_PhiAck/phi_stmt_1690_ack
      -- 
    phi_stmt_1690_ack_12291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 931_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1690_ack_0, ack => minSumDecode_CP_6680_elements(931)); -- 
    -- CP-element group 932:  fork  transition  output  bypass 
    -- CP-element group 932: predecessors 
    -- CP-element group 932: 	24 
    -- CP-element group 932: successors 
    -- CP-element group 932: 	933 
    -- CP-element group 932: 	935 
    -- CP-element group 932: 	936 
    -- CP-element group 932: 	938 
    -- CP-element group 932: 	939 
    -- CP-element group 932:  members (19) 
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Sample/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Sample/rr
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Update/cr
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Sample/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Sample/rr
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Update/cr
      -- 
    rr_12318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(932), ack => type_cast_1712_inst_req_0); -- 
    cr_12323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(932), ack => type_cast_1712_inst_req_1); -- 
    rr_12341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(932), ack => type_cast_1718_inst_req_0); -- 
    cr_12346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(932), ack => type_cast_1718_inst_req_1); -- 
    minSumDecode_CP_6680_elements(932) <= minSumDecode_CP_6680_elements(24);
    -- CP-element group 933:  transition  bypass 
    -- CP-element group 933: predecessors 
    -- CP-element group 933: 	932 
    -- CP-element group 933: successors 
    -- CP-element group 933: 	934 
    -- CP-element group 933:  members (1) 
      -- CP-element group 933: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1704_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(933) is a control-delay.
    cp_element_933_delay: control_delay_element  generic map(name => " 933_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(932), ack => minSumDecode_CP_6680_elements(933), clk => clk, reset =>reset);
    -- CP-element group 934:  transition  output  bypass 
    -- CP-element group 934: predecessors 
    -- CP-element group 934: 	933 
    -- CP-element group 934: successors 
    -- CP-element group 934: 	941 
    -- CP-element group 934:  members (3) 
      -- CP-element group 934: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/$exit
      -- CP-element group 934: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/$exit
      -- CP-element group 934: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_req
      -- 
    phi_stmt_1700_req_12302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1700_req_12302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(934), ack => phi_stmt_1700_req_0); -- 
    minSumDecode_CP_6680_elements(934) <= minSumDecode_CP_6680_elements(933);
    -- CP-element group 935:  transition  input  no-bypass 
    -- CP-element group 935: predecessors 
    -- CP-element group 935: 	932 
    -- CP-element group 935: successors 
    -- CP-element group 935: 	937 
    -- CP-element group 935:  members (2) 
      -- CP-element group 935: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Sample/$exit
      -- CP-element group 935: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Sample/ra
      -- 
    ra_12319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 935_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1712_inst_ack_0, ack => minSumDecode_CP_6680_elements(935)); -- 
    -- CP-element group 936:  transition  input  no-bypass 
    -- CP-element group 936: predecessors 
    -- CP-element group 936: 	932 
    -- CP-element group 936: successors 
    -- CP-element group 936: 	937 
    -- CP-element group 936:  members (2) 
      -- CP-element group 936: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Update/$exit
      -- CP-element group 936: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/Update/ca
      -- 
    ca_12324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 936_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1712_inst_ack_1, ack => minSumDecode_CP_6680_elements(936)); -- 
    -- CP-element group 937:  join  transition  output  bypass 
    -- CP-element group 937: predecessors 
    -- CP-element group 937: 	935 
    -- CP-element group 937: 	936 
    -- CP-element group 937: successors 
    -- CP-element group 937: 	941 
    -- CP-element group 937:  members (5) 
      -- CP-element group 937: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/$exit
      -- CP-element group 937: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$exit
      -- CP-element group 937: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/$exit
      -- CP-element group 937: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1712/SplitProtocol/$exit
      -- CP-element group 937: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_req
      -- 
    phi_stmt_1707_req_12325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1707_req_12325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(937), ack => phi_stmt_1707_req_1); -- 
    minSumDecode_cp_element_group_937: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_937"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(935) & minSumDecode_CP_6680_elements(936);
      gj_minSumDecode_cp_element_group_937 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(937), clk => clk, reset => reset); --
    end block;
    -- CP-element group 938:  transition  input  no-bypass 
    -- CP-element group 938: predecessors 
    -- CP-element group 938: 	932 
    -- CP-element group 938: successors 
    -- CP-element group 938: 	940 
    -- CP-element group 938:  members (2) 
      -- CP-element group 938: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Sample/$exit
      -- CP-element group 938: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Sample/ra
      -- 
    ra_12342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 938_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_0, ack => minSumDecode_CP_6680_elements(938)); -- 
    -- CP-element group 939:  transition  input  no-bypass 
    -- CP-element group 939: predecessors 
    -- CP-element group 939: 	932 
    -- CP-element group 939: successors 
    -- CP-element group 939: 	940 
    -- CP-element group 939:  members (2) 
      -- CP-element group 939: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Update/$exit
      -- CP-element group 939: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/Update/ca
      -- 
    ca_12347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 939_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_1, ack => minSumDecode_CP_6680_elements(939)); -- 
    -- CP-element group 940:  join  transition  output  bypass 
    -- CP-element group 940: predecessors 
    -- CP-element group 940: 	938 
    -- CP-element group 940: 	939 
    -- CP-element group 940: successors 
    -- CP-element group 940: 	941 
    -- CP-element group 940:  members (5) 
      -- CP-element group 940: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/$exit
      -- CP-element group 940: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/$exit
      -- CP-element group 940: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/$exit
      -- CP-element group 940: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1718/SplitProtocol/$exit
      -- CP-element group 940: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_req
      -- 
    phi_stmt_1713_req_12348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1713_req_12348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(940), ack => phi_stmt_1713_req_1); -- 
    minSumDecode_cp_element_group_940: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_940"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(938) & minSumDecode_CP_6680_elements(939);
      gj_minSumDecode_cp_element_group_940 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(940), clk => clk, reset => reset); --
    end block;
    -- CP-element group 941:  join  transition  no-bypass 
    -- CP-element group 941: predecessors 
    -- CP-element group 941: 	934 
    -- CP-element group 941: 	937 
    -- CP-element group 941: 	940 
    -- CP-element group 941: successors 
    -- CP-element group 941: 	953 
    -- CP-element group 941:  members (1) 
      -- CP-element group 941: 	 branch_block_stmt_1353/initializeMessagex_xexitx_xpreheader_initializeMessagex_xexit_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_941: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_941"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(934) & minSumDecode_CP_6680_elements(937) & minSumDecode_CP_6680_elements(940);
      gj_minSumDecode_cp_element_group_941 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(941), clk => clk, reset => reset); --
    end block;
    -- CP-element group 942:  fork  transition  output  bypass 
    -- CP-element group 942: predecessors 
    -- CP-element group 942: 	96 
    -- CP-element group 942: successors 
    -- CP-element group 942: 	943 
    -- CP-element group 942: 	944 
    -- CP-element group 942: 	946 
    -- CP-element group 942: 	947 
    -- CP-element group 942: 	949 
    -- CP-element group 942: 	950 
    -- CP-element group 942:  members (25) 
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Sample/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Sample/rr
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Update/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Update/cr
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/rr
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/cr
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Sample/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Sample/rr
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Update/$entry
      -- CP-element group 942: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Update/cr
      -- 
    rr_12367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1706_inst_req_0); -- 
    cr_12372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1706_inst_req_1); -- 
    rr_12390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1710_inst_req_0); -- 
    cr_12395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1710_inst_req_1); -- 
    rr_12413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1716_inst_req_0); -- 
    cr_12418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(942), ack => type_cast_1716_inst_req_1); -- 
    minSumDecode_CP_6680_elements(942) <= minSumDecode_CP_6680_elements(96);
    -- CP-element group 943:  transition  input  no-bypass 
    -- CP-element group 943: predecessors 
    -- CP-element group 943: 	942 
    -- CP-element group 943: successors 
    -- CP-element group 943: 	945 
    -- CP-element group 943:  members (2) 
      -- CP-element group 943: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Sample/$exit
      -- CP-element group 943: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Sample/ra
      -- 
    ra_12368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 943_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_0, ack => minSumDecode_CP_6680_elements(943)); -- 
    -- CP-element group 944:  transition  input  no-bypass 
    -- CP-element group 944: predecessors 
    -- CP-element group 944: 	942 
    -- CP-element group 944: successors 
    -- CP-element group 944: 	945 
    -- CP-element group 944:  members (2) 
      -- CP-element group 944: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Update/$exit
      -- CP-element group 944: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/Update/ca
      -- 
    ca_12373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 944_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_1, ack => minSumDecode_CP_6680_elements(944)); -- 
    -- CP-element group 945:  join  transition  output  bypass 
    -- CP-element group 945: predecessors 
    -- CP-element group 945: 	943 
    -- CP-element group 945: 	944 
    -- CP-element group 945: successors 
    -- CP-element group 945: 	952 
    -- CP-element group 945:  members (5) 
      -- CP-element group 945: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/$exit
      -- CP-element group 945: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/$exit
      -- CP-element group 945: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/$exit
      -- CP-element group 945: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_sources/type_cast_1706/SplitProtocol/$exit
      -- CP-element group 945: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1700/phi_stmt_1700_req
      -- 
    phi_stmt_1700_req_12374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1700_req_12374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(945), ack => phi_stmt_1700_req_1); -- 
    minSumDecode_cp_element_group_945: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_945"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(943) & minSumDecode_CP_6680_elements(944);
      gj_minSumDecode_cp_element_group_945 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(945), clk => clk, reset => reset); --
    end block;
    -- CP-element group 946:  transition  input  no-bypass 
    -- CP-element group 946: predecessors 
    -- CP-element group 946: 	942 
    -- CP-element group 946: successors 
    -- CP-element group 946: 	948 
    -- CP-element group 946:  members (2) 
      -- CP-element group 946: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/$exit
      -- CP-element group 946: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/ra
      -- 
    ra_12391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 946_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_0, ack => minSumDecode_CP_6680_elements(946)); -- 
    -- CP-element group 947:  transition  input  no-bypass 
    -- CP-element group 947: predecessors 
    -- CP-element group 947: 	942 
    -- CP-element group 947: successors 
    -- CP-element group 947: 	948 
    -- CP-element group 947:  members (2) 
      -- CP-element group 947: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/$exit
      -- CP-element group 947: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/ca
      -- 
    ca_12396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 947_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_1, ack => minSumDecode_CP_6680_elements(947)); -- 
    -- CP-element group 948:  join  transition  output  bypass 
    -- CP-element group 948: predecessors 
    -- CP-element group 948: 	946 
    -- CP-element group 948: 	947 
    -- CP-element group 948: successors 
    -- CP-element group 948: 	952 
    -- CP-element group 948:  members (5) 
      -- CP-element group 948: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/$exit
      -- CP-element group 948: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$exit
      -- CP-element group 948: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/$exit
      -- CP-element group 948: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/$exit
      -- CP-element group 948: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1707/phi_stmt_1707_req
      -- 
    phi_stmt_1707_req_12397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1707_req_12397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(948), ack => phi_stmt_1707_req_0); -- 
    minSumDecode_cp_element_group_948: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_948"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(946) & minSumDecode_CP_6680_elements(947);
      gj_minSumDecode_cp_element_group_948 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(948), clk => clk, reset => reset); --
    end block;
    -- CP-element group 949:  transition  input  no-bypass 
    -- CP-element group 949: predecessors 
    -- CP-element group 949: 	942 
    -- CP-element group 949: successors 
    -- CP-element group 949: 	951 
    -- CP-element group 949:  members (2) 
      -- CP-element group 949: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Sample/$exit
      -- CP-element group 949: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Sample/ra
      -- 
    ra_12414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 949_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_0, ack => minSumDecode_CP_6680_elements(949)); -- 
    -- CP-element group 950:  transition  input  no-bypass 
    -- CP-element group 950: predecessors 
    -- CP-element group 950: 	942 
    -- CP-element group 950: successors 
    -- CP-element group 950: 	951 
    -- CP-element group 950:  members (2) 
      -- CP-element group 950: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Update/$exit
      -- CP-element group 950: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/Update/ca
      -- 
    ca_12419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 950_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_1, ack => minSumDecode_CP_6680_elements(950)); -- 
    -- CP-element group 951:  join  transition  output  bypass 
    -- CP-element group 951: predecessors 
    -- CP-element group 951: 	949 
    -- CP-element group 951: 	950 
    -- CP-element group 951: successors 
    -- CP-element group 951: 	952 
    -- CP-element group 951:  members (5) 
      -- CP-element group 951: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/$exit
      -- CP-element group 951: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/$exit
      -- CP-element group 951: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/$exit
      -- CP-element group 951: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_sources/type_cast_1716/SplitProtocol/$exit
      -- CP-element group 951: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/phi_stmt_1713/phi_stmt_1713_req
      -- 
    phi_stmt_1713_req_12420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1713_req_12420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(951), ack => phi_stmt_1713_req_0); -- 
    minSumDecode_cp_element_group_951: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_951"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(949) & minSumDecode_CP_6680_elements(950);
      gj_minSumDecode_cp_element_group_951 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(951), clk => clk, reset => reset); --
    end block;
    -- CP-element group 952:  join  transition  bypass 
    -- CP-element group 952: predecessors 
    -- CP-element group 952: 	945 
    -- CP-element group 952: 	948 
    -- CP-element group 952: 	951 
    -- CP-element group 952: successors 
    -- CP-element group 952: 	953 
    -- CP-element group 952:  members (1) 
      -- CP-element group 952: 	 branch_block_stmt_1353/updateMessagex_xexit_initializeMessagex_xexit_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_952: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_952"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(945) & minSumDecode_CP_6680_elements(948) & minSumDecode_CP_6680_elements(951);
      gj_minSumDecode_cp_element_group_952 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(952), clk => clk, reset => reset); --
    end block;
    -- CP-element group 953:  merge  place  bypass 
    -- CP-element group 953: predecessors 
    -- CP-element group 953: 	941 
    -- CP-element group 953: 	952 
    -- CP-element group 953: successors 
    -- CP-element group 953: 	954 
    -- CP-element group 953:  members (1) 
      -- CP-element group 953: 	 branch_block_stmt_1353/merge_stmt_1699_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(953) <= OrReduce(minSumDecode_CP_6680_elements(941) & minSumDecode_CP_6680_elements(952));
    -- CP-element group 954:  fork  transition  bypass 
    -- CP-element group 954: predecessors 
    -- CP-element group 954: 	953 
    -- CP-element group 954: successors 
    -- CP-element group 954: 	955 
    -- CP-element group 954: 	956 
    -- CP-element group 954: 	957 
    -- CP-element group 954:  members (1) 
      -- CP-element group 954: 	 branch_block_stmt_1353/merge_stmt_1699_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(954) <= minSumDecode_CP_6680_elements(953);
    -- CP-element group 955:  transition  input  no-bypass 
    -- CP-element group 955: predecessors 
    -- CP-element group 955: 	954 
    -- CP-element group 955: successors 
    -- CP-element group 955: 	958 
    -- CP-element group 955:  members (1) 
      -- CP-element group 955: 	 branch_block_stmt_1353/merge_stmt_1699_PhiAck/phi_stmt_1700_ack
      -- 
    phi_stmt_1700_ack_12425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 955_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1700_ack_0, ack => minSumDecode_CP_6680_elements(955)); -- 
    -- CP-element group 956:  transition  input  no-bypass 
    -- CP-element group 956: predecessors 
    -- CP-element group 956: 	954 
    -- CP-element group 956: successors 
    -- CP-element group 956: 	958 
    -- CP-element group 956:  members (1) 
      -- CP-element group 956: 	 branch_block_stmt_1353/merge_stmt_1699_PhiAck/phi_stmt_1707_ack
      -- 
    phi_stmt_1707_ack_12426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 956_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1707_ack_0, ack => minSumDecode_CP_6680_elements(956)); -- 
    -- CP-element group 957:  transition  input  no-bypass 
    -- CP-element group 957: predecessors 
    -- CP-element group 957: 	954 
    -- CP-element group 957: successors 
    -- CP-element group 957: 	958 
    -- CP-element group 957:  members (1) 
      -- CP-element group 957: 	 branch_block_stmt_1353/merge_stmt_1699_PhiAck/phi_stmt_1713_ack
      -- 
    phi_stmt_1713_ack_12427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 957_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1713_ack_0, ack => minSumDecode_CP_6680_elements(957)); -- 
    -- CP-element group 958:  join  transition  bypass 
    -- CP-element group 958: predecessors 
    -- CP-element group 958: 	955 
    -- CP-element group 958: 	956 
    -- CP-element group 958: 	957 
    -- CP-element group 958: successors 
    -- CP-element group 958: 	25 
    -- CP-element group 958:  members (1) 
      -- CP-element group 958: 	 branch_block_stmt_1353/merge_stmt_1699_PhiAck/$exit
      -- 
    minSumDecode_cp_element_group_958: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_958"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(955) & minSumDecode_CP_6680_elements(956) & minSumDecode_CP_6680_elements(957);
      gj_minSumDecode_cp_element_group_958 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(958), clk => clk, reset => reset); --
    end block;
    -- CP-element group 959:  transition  bypass 
    -- CP-element group 959: predecessors 
    -- CP-element group 959: 	351 
    -- CP-element group 959: successors 
    -- CP-element group 959: 	960 
    -- CP-element group 959:  members (2) 
      -- CP-element group 959: 	 branch_block_stmt_1353/initializeMessagex_xexit_bb_14_PhiReq/$entry
      -- CP-element group 959: 	 branch_block_stmt_1353/initializeMessagex_xexit_bb_14_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(959) <= minSumDecode_CP_6680_elements(351);
    -- CP-element group 960:  place  bypass 
    -- CP-element group 960: predecessors 
    -- CP-element group 960: 	959 
    -- CP-element group 960: successors 
    -- CP-element group 960: 	961 
    -- CP-element group 960:  members (1) 
      -- CP-element group 960: 	 branch_block_stmt_1353/merge_stmt_1740_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(960) <= minSumDecode_CP_6680_elements(959);
    -- CP-element group 961:  transition  bypass 
    -- CP-element group 961: predecessors 
    -- CP-element group 961: 	960 
    -- CP-element group 961: successors 
    -- CP-element group 961: 	27 
    -- CP-element group 961:  members (3) 
      -- CP-element group 961: 	 branch_block_stmt_1353/merge_stmt_1740_PhiAck/$entry
      -- CP-element group 961: 	 branch_block_stmt_1353/merge_stmt_1740_PhiAck/$exit
      -- CP-element group 961: 	 branch_block_stmt_1353/merge_stmt_1740_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(961) <= minSumDecode_CP_6680_elements(960);
    -- CP-element group 962:  transition  bypass 
    -- CP-element group 962: predecessors 
    -- CP-element group 962: 	364 
    -- CP-element group 962: successors 
    -- CP-element group 962: 	963 
    -- CP-element group 962:  members (2) 
      -- CP-element group 962: 	 branch_block_stmt_1353/bb_14_bbx_xnphx_xi18_PhiReq/$entry
      -- CP-element group 962: 	 branch_block_stmt_1353/bb_14_bbx_xnphx_xi18_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(962) <= minSumDecode_CP_6680_elements(364);
    -- CP-element group 963:  place  bypass 
    -- CP-element group 963: predecessors 
    -- CP-element group 963: 	962 
    -- CP-element group 963: successors 
    -- CP-element group 963: 	964 
    -- CP-element group 963:  members (1) 
      -- CP-element group 963: 	 branch_block_stmt_1353/merge_stmt_1753_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(963) <= minSumDecode_CP_6680_elements(962);
    -- CP-element group 964:  transition  bypass 
    -- CP-element group 964: predecessors 
    -- CP-element group 964: 	963 
    -- CP-element group 964: successors 
    -- CP-element group 964: 	29 
    -- CP-element group 964:  members (3) 
      -- CP-element group 964: 	 branch_block_stmt_1353/merge_stmt_1753_PhiAck/$entry
      -- CP-element group 964: 	 branch_block_stmt_1353/merge_stmt_1753_PhiAck/$exit
      -- CP-element group 964: 	 branch_block_stmt_1353/merge_stmt_1753_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(964) <= minSumDecode_CP_6680_elements(963);
    -- CP-element group 965:  fork  transition  output  bypass 
    -- CP-element group 965: predecessors 
    -- CP-element group 965: 	401 
    -- CP-element group 965: successors 
    -- CP-element group 965: 	966 
    -- CP-element group 965: 	967 
    -- CP-element group 965:  members (9) 
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Sample/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Sample/rr
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Update/$entry
      -- CP-element group 965: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Update/cr
      -- 
    rr_12470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(965), ack => type_cast_1791_inst_req_0); -- 
    cr_12475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(965), ack => type_cast_1791_inst_req_1); -- 
    minSumDecode_CP_6680_elements(965) <= minSumDecode_CP_6680_elements(401);
    -- CP-element group 966:  transition  input  no-bypass 
    -- CP-element group 966: predecessors 
    -- CP-element group 966: 	965 
    -- CP-element group 966: successors 
    -- CP-element group 966: 	968 
    -- CP-element group 966:  members (2) 
      -- CP-element group 966: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Sample/$exit
      -- CP-element group 966: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Sample/ra
      -- 
    ra_12471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 966_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_0, ack => minSumDecode_CP_6680_elements(966)); -- 
    -- CP-element group 967:  transition  input  no-bypass 
    -- CP-element group 967: predecessors 
    -- CP-element group 967: 	965 
    -- CP-element group 967: successors 
    -- CP-element group 967: 	968 
    -- CP-element group 967:  members (2) 
      -- CP-element group 967: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Update/$exit
      -- CP-element group 967: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/Update/ca
      -- 
    ca_12476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 967_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_1, ack => minSumDecode_CP_6680_elements(967)); -- 
    -- CP-element group 968:  join  transition  output  bypass 
    -- CP-element group 968: predecessors 
    -- CP-element group 968: 	966 
    -- CP-element group 968: 	967 
    -- CP-element group 968: successors 
    -- CP-element group 968: 	972 
    -- CP-element group 968:  members (6) 
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/$exit
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/$exit
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/$exit
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/$exit
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1791/SplitProtocol/$exit
      -- CP-element group 968: 	 branch_block_stmt_1353/bb_16_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_req
      -- 
    phi_stmt_1785_req_12477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1785_req_12477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(968), ack => phi_stmt_1785_req_1); -- 
    minSumDecode_cp_element_group_968: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_968"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(966) & minSumDecode_CP_6680_elements(967);
      gj_minSumDecode_cp_element_group_968 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(968), clk => clk, reset => reset); --
    end block;
    -- CP-element group 969:  transition  bypass 
    -- CP-element group 969: predecessors 
    -- CP-element group 969: 	30 
    -- CP-element group 969: successors 
    -- CP-element group 969: 	970 
    -- CP-element group 969:  members (3) 
      -- CP-element group 969: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/$entry
      -- CP-element group 969: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/$entry
      -- CP-element group 969: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(969) <= minSumDecode_CP_6680_elements(30);
    -- CP-element group 970:  transition  bypass 
    -- CP-element group 970: predecessors 
    -- CP-element group 970: 	969 
    -- CP-element group 970: successors 
    -- CP-element group 970: 	971 
    -- CP-element group 970:  members (1) 
      -- CP-element group 970: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/type_cast_1789_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(970) is a control-delay.
    cp_element_970_delay: control_delay_element  generic map(name => " 970_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(969), ack => minSumDecode_CP_6680_elements(970), clk => clk, reset =>reset);
    -- CP-element group 971:  transition  output  bypass 
    -- CP-element group 971: predecessors 
    -- CP-element group 971: 	970 
    -- CP-element group 971: successors 
    -- CP-element group 971: 	972 
    -- CP-element group 971:  members (4) 
      -- CP-element group 971: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/$exit
      -- CP-element group 971: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/$exit
      -- CP-element group 971: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_sources/$exit
      -- CP-element group 971: 	 branch_block_stmt_1353/bbx_xnphx_xi18_bb_16_PhiReq/phi_stmt_1785/phi_stmt_1785_req
      -- 
    phi_stmt_1785_req_12488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1785_req_12488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(971), ack => phi_stmt_1785_req_0); -- 
    minSumDecode_CP_6680_elements(971) <= minSumDecode_CP_6680_elements(970);
    -- CP-element group 972:  merge  place  bypass 
    -- CP-element group 972: predecessors 
    -- CP-element group 972: 	968 
    -- CP-element group 972: 	971 
    -- CP-element group 972: successors 
    -- CP-element group 972: 	973 
    -- CP-element group 972:  members (1) 
      -- CP-element group 972: 	 branch_block_stmt_1353/merge_stmt_1784_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(972) <= OrReduce(minSumDecode_CP_6680_elements(968) & minSumDecode_CP_6680_elements(971));
    -- CP-element group 973:  transition  bypass 
    -- CP-element group 973: predecessors 
    -- CP-element group 973: 	972 
    -- CP-element group 973: successors 
    -- CP-element group 973: 	974 
    -- CP-element group 973:  members (1) 
      -- CP-element group 973: 	 branch_block_stmt_1353/merge_stmt_1784_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(973) <= minSumDecode_CP_6680_elements(972);
    -- CP-element group 974:  transition  input  no-bypass 
    -- CP-element group 974: predecessors 
    -- CP-element group 974: 	973 
    -- CP-element group 974: successors 
    -- CP-element group 974: 	31 
    -- CP-element group 974:  members (2) 
      -- CP-element group 974: 	 branch_block_stmt_1353/merge_stmt_1784_PhiAck/$exit
      -- CP-element group 974: 	 branch_block_stmt_1353/merge_stmt_1784_PhiAck/phi_stmt_1785_ack
      -- 
    phi_stmt_1785_ack_12493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 974_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1785_ack_0, ack => minSumDecode_CP_6680_elements(974)); -- 
    -- CP-element group 975:  transition  bypass 
    -- CP-element group 975: predecessors 
    -- CP-element group 975: 	400 
    -- CP-element group 975: successors 
    -- CP-element group 975: 	976 
    -- CP-element group 975:  members (2) 
      -- CP-element group 975: 	 branch_block_stmt_1353/bb_16_initialize_aPosteriorix_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 975: 	 branch_block_stmt_1353/bb_16_initialize_aPosteriorix_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(975) <= minSumDecode_CP_6680_elements(400);
    -- CP-element group 976:  place  bypass 
    -- CP-element group 976: predecessors 
    -- CP-element group 976: 	975 
    -- CP-element group 976: successors 
    -- CP-element group 976: 	977 
    -- CP-element group 976:  members (1) 
      -- CP-element group 976: 	 branch_block_stmt_1353/merge_stmt_1828_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(976) <= minSumDecode_CP_6680_elements(975);
    -- CP-element group 977:  transition  bypass 
    -- CP-element group 977: predecessors 
    -- CP-element group 977: 	976 
    -- CP-element group 977: successors 
    -- CP-element group 977: 	33 
    -- CP-element group 977:  members (3) 
      -- CP-element group 977: 	 branch_block_stmt_1353/merge_stmt_1828_PhiAck/$entry
      -- CP-element group 977: 	 branch_block_stmt_1353/merge_stmt_1828_PhiAck/$exit
      -- CP-element group 977: 	 branch_block_stmt_1353/merge_stmt_1828_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(977) <= minSumDecode_CP_6680_elements(976);
    -- CP-element group 978:  transition  bypass 
    -- CP-element group 978: predecessors 
    -- CP-element group 978: 	363 
    -- CP-element group 978: successors 
    -- CP-element group 978: 	980 
    -- CP-element group 978:  members (2) 
      -- CP-element group 978: 	 branch_block_stmt_1353/bb_14_initialize_aPosteriorix_xexit_PhiReq/$entry
      -- CP-element group 978: 	 branch_block_stmt_1353/bb_14_initialize_aPosteriorix_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(978) <= minSumDecode_CP_6680_elements(363);
    -- CP-element group 979:  transition  bypass 
    -- CP-element group 979: predecessors 
    -- CP-element group 979: 	33 
    -- CP-element group 979: successors 
    -- CP-element group 979: 	980 
    -- CP-element group 979:  members (2) 
      -- CP-element group 979: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexitx_xloopexit_initialize_aPosteriorix_xexit_PhiReq/$entry
      -- CP-element group 979: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexitx_xloopexit_initialize_aPosteriorix_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(979) <= minSumDecode_CP_6680_elements(33);
    -- CP-element group 980:  merge  place  bypass 
    -- CP-element group 980: predecessors 
    -- CP-element group 980: 	978 
    -- CP-element group 980: 	979 
    -- CP-element group 980: successors 
    -- CP-element group 980: 	981 
    -- CP-element group 980:  members (1) 
      -- CP-element group 980: 	 branch_block_stmt_1353/merge_stmt_1830_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(980) <= OrReduce(minSumDecode_CP_6680_elements(978) & minSumDecode_CP_6680_elements(979));
    -- CP-element group 981:  transition  bypass 
    -- CP-element group 981: predecessors 
    -- CP-element group 981: 	980 
    -- CP-element group 981: successors 
    -- CP-element group 981: 	34 
    -- CP-element group 981:  members (3) 
      -- CP-element group 981: 	 branch_block_stmt_1353/merge_stmt_1830_PhiAck/$entry
      -- CP-element group 981: 	 branch_block_stmt_1353/merge_stmt_1830_PhiAck/$exit
      -- CP-element group 981: 	 branch_block_stmt_1353/merge_stmt_1830_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(981) <= minSumDecode_CP_6680_elements(980);
    -- CP-element group 982:  transition  bypass 
    -- CP-element group 982: predecessors 
    -- CP-element group 982: 	413 
    -- CP-element group 982: successors 
    -- CP-element group 982: 	983 
    -- CP-element group 982:  members (2) 
      -- CP-element group 982: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_bbx_xnphx_xi27_PhiReq/$entry
      -- CP-element group 982: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_bbx_xnphx_xi27_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(982) <= minSumDecode_CP_6680_elements(413);
    -- CP-element group 983:  place  bypass 
    -- CP-element group 983: predecessors 
    -- CP-element group 983: 	982 
    -- CP-element group 983: successors 
    -- CP-element group 983: 	984 
    -- CP-element group 983:  members (1) 
      -- CP-element group 983: 	 branch_block_stmt_1353/merge_stmt_1843_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(983) <= minSumDecode_CP_6680_elements(982);
    -- CP-element group 984:  transition  bypass 
    -- CP-element group 984: predecessors 
    -- CP-element group 984: 	983 
    -- CP-element group 984: successors 
    -- CP-element group 984: 	36 
    -- CP-element group 984:  members (3) 
      -- CP-element group 984: 	 branch_block_stmt_1353/merge_stmt_1843_PhiAck/$entry
      -- CP-element group 984: 	 branch_block_stmt_1353/merge_stmt_1843_PhiAck/$exit
      -- CP-element group 984: 	 branch_block_stmt_1353/merge_stmt_1843_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(984) <= minSumDecode_CP_6680_elements(983);
    -- CP-element group 985:  fork  transition  output  bypass 
    -- CP-element group 985: predecessors 
    -- CP-element group 985: 	445 
    -- CP-element group 985: successors 
    -- CP-element group 985: 	986 
    -- CP-element group 985: 	987 
    -- CP-element group 985:  members (9) 
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/rr
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/$entry
      -- CP-element group 985: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/cr
      -- 
    rr_12547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(985), ack => type_cast_1881_inst_req_0); -- 
    cr_12552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(985), ack => type_cast_1881_inst_req_1); -- 
    minSumDecode_CP_6680_elements(985) <= minSumDecode_CP_6680_elements(445);
    -- CP-element group 986:  transition  input  no-bypass 
    -- CP-element group 986: predecessors 
    -- CP-element group 986: 	985 
    -- CP-element group 986: successors 
    -- CP-element group 986: 	988 
    -- CP-element group 986:  members (2) 
      -- CP-element group 986: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/$exit
      -- CP-element group 986: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/ra
      -- 
    ra_12548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 986_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_0, ack => minSumDecode_CP_6680_elements(986)); -- 
    -- CP-element group 987:  transition  input  no-bypass 
    -- CP-element group 987: predecessors 
    -- CP-element group 987: 	985 
    -- CP-element group 987: successors 
    -- CP-element group 987: 	988 
    -- CP-element group 987:  members (2) 
      -- CP-element group 987: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/$exit
      -- CP-element group 987: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/ca
      -- 
    ca_12553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 987_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_1, ack => minSumDecode_CP_6680_elements(987)); -- 
    -- CP-element group 988:  join  transition  output  bypass 
    -- CP-element group 988: predecessors 
    -- CP-element group 988: 	986 
    -- CP-element group 988: 	987 
    -- CP-element group 988: successors 
    -- CP-element group 988: 	992 
    -- CP-element group 988:  members (6) 
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/$exit
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/$exit
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/$exit
      -- CP-element group 988: 	 branch_block_stmt_1353/bb_20_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_12554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_12554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(988), ack => phi_stmt_1875_req_1); -- 
    minSumDecode_cp_element_group_988: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "minSumDecode_cp_element_group_988"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(986) & minSumDecode_CP_6680_elements(987);
      gj_minSumDecode_cp_element_group_988 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(988), clk => clk, reset => reset); --
    end block;
    -- CP-element group 989:  transition  bypass 
    -- CP-element group 989: predecessors 
    -- CP-element group 989: 	37 
    -- CP-element group 989: successors 
    -- CP-element group 989: 	990 
    -- CP-element group 989:  members (3) 
      -- CP-element group 989: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/$entry
      -- CP-element group 989: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 989: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(989) <= minSumDecode_CP_6680_elements(37);
    -- CP-element group 990:  transition  bypass 
    -- CP-element group 990: predecessors 
    -- CP-element group 990: 	989 
    -- CP-element group 990: successors 
    -- CP-element group 990: 	991 
    -- CP-element group 990:  members (1) 
      -- CP-element group 990: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1879_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(990) is a control-delay.
    cp_element_990_delay: control_delay_element  generic map(name => " 990_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(989), ack => minSumDecode_CP_6680_elements(990), clk => clk, reset =>reset);
    -- CP-element group 991:  transition  output  bypass 
    -- CP-element group 991: predecessors 
    -- CP-element group 991: 	990 
    -- CP-element group 991: successors 
    -- CP-element group 991: 	992 
    -- CP-element group 991:  members (4) 
      -- CP-element group 991: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/$exit
      -- CP-element group 991: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 991: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 991: 	 branch_block_stmt_1353/bbx_xnphx_xi27_bb_20_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_12565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_12565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(991), ack => phi_stmt_1875_req_0); -- 
    minSumDecode_CP_6680_elements(991) <= minSumDecode_CP_6680_elements(990);
    -- CP-element group 992:  merge  place  bypass 
    -- CP-element group 992: predecessors 
    -- CP-element group 992: 	988 
    -- CP-element group 992: 	991 
    -- CP-element group 992: successors 
    -- CP-element group 992: 	993 
    -- CP-element group 992:  members (1) 
      -- CP-element group 992: 	 branch_block_stmt_1353/merge_stmt_1874_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(992) <= OrReduce(minSumDecode_CP_6680_elements(988) & minSumDecode_CP_6680_elements(991));
    -- CP-element group 993:  transition  bypass 
    -- CP-element group 993: predecessors 
    -- CP-element group 993: 	992 
    -- CP-element group 993: successors 
    -- CP-element group 993: 	994 
    -- CP-element group 993:  members (1) 
      -- CP-element group 993: 	 branch_block_stmt_1353/merge_stmt_1874_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(993) <= minSumDecode_CP_6680_elements(992);
    -- CP-element group 994:  transition  input  no-bypass 
    -- CP-element group 994: predecessors 
    -- CP-element group 994: 	993 
    -- CP-element group 994: successors 
    -- CP-element group 994: 	38 
    -- CP-element group 994:  members (2) 
      -- CP-element group 994: 	 branch_block_stmt_1353/merge_stmt_1874_PhiAck/$exit
      -- CP-element group 994: 	 branch_block_stmt_1353/merge_stmt_1874_PhiAck/phi_stmt_1875_ack
      -- 
    phi_stmt_1875_ack_12570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 994_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1875_ack_0, ack => minSumDecode_CP_6680_elements(994)); -- 
    -- CP-element group 995:  transition  bypass 
    -- CP-element group 995: predecessors 
    -- CP-element group 995: 	444 
    -- CP-element group 995: successors 
    -- CP-element group 995: 	996 
    -- CP-element group 995:  members (2) 
      -- CP-element group 995: 	 branch_block_stmt_1353/bb_20_initializeExtrinsicInfox_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 995: 	 branch_block_stmt_1353/bb_20_initializeExtrinsicInfox_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(995) <= minSumDecode_CP_6680_elements(444);
    -- CP-element group 996:  place  bypass 
    -- CP-element group 996: predecessors 
    -- CP-element group 996: 	995 
    -- CP-element group 996: successors 
    -- CP-element group 996: 	997 
    -- CP-element group 996:  members (1) 
      -- CP-element group 996: 	 branch_block_stmt_1353/merge_stmt_1910_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(996) <= minSumDecode_CP_6680_elements(995);
    -- CP-element group 997:  transition  bypass 
    -- CP-element group 997: predecessors 
    -- CP-element group 997: 	996 
    -- CP-element group 997: successors 
    -- CP-element group 997: 	40 
    -- CP-element group 997:  members (3) 
      -- CP-element group 997: 	 branch_block_stmt_1353/merge_stmt_1910_PhiAck/$entry
      -- CP-element group 997: 	 branch_block_stmt_1353/merge_stmt_1910_PhiAck/$exit
      -- CP-element group 997: 	 branch_block_stmt_1353/merge_stmt_1910_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(997) <= minSumDecode_CP_6680_elements(996);
    -- CP-element group 998:  transition  bypass 
    -- CP-element group 998: predecessors 
    -- CP-element group 998: 	40 
    -- CP-element group 998: successors 
    -- CP-element group 998: 	1000 
    -- CP-element group 998:  members (2) 
      -- CP-element group 998: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexitx_xloopexit_initializeExtrinsicInfox_xexit_PhiReq/$entry
      -- CP-element group 998: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexitx_xloopexit_initializeExtrinsicInfox_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(998) <= minSumDecode_CP_6680_elements(40);
    -- CP-element group 999:  transition  bypass 
    -- CP-element group 999: predecessors 
    -- CP-element group 999: 	412 
    -- CP-element group 999: successors 
    -- CP-element group 999: 	1000 
    -- CP-element group 999:  members (2) 
      -- CP-element group 999: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_initializeExtrinsicInfox_xexit_PhiReq/$entry
      -- CP-element group 999: 	 branch_block_stmt_1353/initialize_aPosteriorix_xexit_initializeExtrinsicInfox_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(999) <= minSumDecode_CP_6680_elements(412);
    -- CP-element group 1000:  merge  place  bypass 
    -- CP-element group 1000: predecessors 
    -- CP-element group 1000: 	998 
    -- CP-element group 1000: 	999 
    -- CP-element group 1000: successors 
    -- CP-element group 1000: 	1001 
    -- CP-element group 1000:  members (1) 
      -- CP-element group 1000: 	 branch_block_stmt_1353/merge_stmt_1912_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1000) <= OrReduce(minSumDecode_CP_6680_elements(998) & minSumDecode_CP_6680_elements(999));
    -- CP-element group 1001:  transition  bypass 
    -- CP-element group 1001: predecessors 
    -- CP-element group 1001: 	1000 
    -- CP-element group 1001: successors 
    -- CP-element group 1001: 	41 
    -- CP-element group 1001:  members (3) 
      -- CP-element group 1001: 	 branch_block_stmt_1353/merge_stmt_1912_PhiAck/$entry
      -- CP-element group 1001: 	 branch_block_stmt_1353/merge_stmt_1912_PhiAck/$exit
      -- CP-element group 1001: 	 branch_block_stmt_1353/merge_stmt_1912_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1001) <= minSumDecode_CP_6680_elements(1000);
    -- CP-element group 1002:  transition  bypass 
    -- CP-element group 1002: predecessors 
    -- CP-element group 1002: 	462 
    -- CP-element group 1002: successors 
    -- CP-element group 1002: 	1003 
    -- CP-element group 1002:  members (2) 
      -- CP-element group 1002: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_bbx_xnphx_xi54_PhiReq/$entry
      -- CP-element group 1002: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_bbx_xnphx_xi54_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1002) <= minSumDecode_CP_6680_elements(462);
    -- CP-element group 1003:  place  bypass 
    -- CP-element group 1003: predecessors 
    -- CP-element group 1003: 	1002 
    -- CP-element group 1003: successors 
    -- CP-element group 1003: 	1004 
    -- CP-element group 1003:  members (1) 
      -- CP-element group 1003: 	 branch_block_stmt_1353/merge_stmt_1929_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1003) <= minSumDecode_CP_6680_elements(1002);
    -- CP-element group 1004:  transition  bypass 
    -- CP-element group 1004: predecessors 
    -- CP-element group 1004: 	1003 
    -- CP-element group 1004: successors 
    -- CP-element group 1004: 	44 
    -- CP-element group 1004:  members (3) 
      -- CP-element group 1004: 	 branch_block_stmt_1353/merge_stmt_1929_PhiAck/$entry
      -- CP-element group 1004: 	 branch_block_stmt_1353/merge_stmt_1929_PhiAck/$exit
      -- CP-element group 1004: 	 branch_block_stmt_1353/merge_stmt_1929_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1004) <= minSumDecode_CP_6680_elements(1003);
    -- CP-element group 1005:  fork  transition  output  bypass 
    -- CP-element group 1005: predecessors 
    -- CP-element group 1005: 	515 
    -- CP-element group 1005: successors 
    -- CP-element group 1005: 	1006 
    -- CP-element group 1005: 	1007 
    -- CP-element group 1005:  members (9) 
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Sample/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Sample/rr
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Update/$entry
      -- CP-element group 1005: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Update/cr
      -- 
    rr_12624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1005), ack => type_cast_1967_inst_req_0); -- 
    cr_12629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1005), ack => type_cast_1967_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1005) <= minSumDecode_CP_6680_elements(515);
    -- CP-element group 1006:  transition  input  no-bypass 
    -- CP-element group 1006: predecessors 
    -- CP-element group 1006: 	1005 
    -- CP-element group 1006: successors 
    -- CP-element group 1006: 	1008 
    -- CP-element group 1006:  members (2) 
      -- CP-element group 1006: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Sample/$exit
      -- CP-element group 1006: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Sample/ra
      -- 
    ra_12625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1006_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1967_inst_ack_0, ack => minSumDecode_CP_6680_elements(1006)); -- 
    -- CP-element group 1007:  transition  input  no-bypass 
    -- CP-element group 1007: predecessors 
    -- CP-element group 1007: 	1005 
    -- CP-element group 1007: successors 
    -- CP-element group 1007: 	1008 
    -- CP-element group 1007:  members (2) 
      -- CP-element group 1007: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Update/$exit
      -- CP-element group 1007: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/Update/ca
      -- 
    ca_12630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1007_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1967_inst_ack_1, ack => minSumDecode_CP_6680_elements(1007)); -- 
    -- CP-element group 1008:  join  transition  output  bypass 
    -- CP-element group 1008: predecessors 
    -- CP-element group 1008: 	1006 
    -- CP-element group 1008: 	1007 
    -- CP-element group 1008: successors 
    -- CP-element group 1008: 	1012 
    -- CP-element group 1008:  members (6) 
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/$exit
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/$exit
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$exit
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/$exit
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967/SplitProtocol/$exit
      -- CP-element group 1008: 	 branch_block_stmt_1353/bb_24_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_req
      -- 
    phi_stmt_1961_req_12631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1961_req_12631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1008), ack => phi_stmt_1961_req_1); -- 
    minSumDecode_cp_element_group_1008: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1008"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1006) & minSumDecode_CP_6680_elements(1007);
      gj_minSumDecode_cp_element_group_1008 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1008), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1009:  transition  bypass 
    -- CP-element group 1009: predecessors 
    -- CP-element group 1009: 	45 
    -- CP-element group 1009: successors 
    -- CP-element group 1009: 	1010 
    -- CP-element group 1009:  members (3) 
      -- CP-element group 1009: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/$entry
      -- CP-element group 1009: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/$entry
      -- CP-element group 1009: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1009) <= minSumDecode_CP_6680_elements(45);
    -- CP-element group 1010:  transition  bypass 
    -- CP-element group 1010: predecessors 
    -- CP-element group 1010: 	1009 
    -- CP-element group 1010: successors 
    -- CP-element group 1010: 	1011 
    -- CP-element group 1010:  members (1) 
      -- CP-element group 1010: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1965_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1010) is a control-delay.
    cp_element_1010_delay: control_delay_element  generic map(name => " 1010_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1009), ack => minSumDecode_CP_6680_elements(1010), clk => clk, reset =>reset);
    -- CP-element group 1011:  transition  output  bypass 
    -- CP-element group 1011: predecessors 
    -- CP-element group 1011: 	1010 
    -- CP-element group 1011: successors 
    -- CP-element group 1011: 	1012 
    -- CP-element group 1011:  members (4) 
      -- CP-element group 1011: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/$exit
      -- CP-element group 1011: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/$exit
      -- CP-element group 1011: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$exit
      -- CP-element group 1011: 	 branch_block_stmt_1353/bbx_xnphx_xi54_bb_24_PhiReq/phi_stmt_1961/phi_stmt_1961_req
      -- 
    phi_stmt_1961_req_12642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1961_req_12642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1011), ack => phi_stmt_1961_req_0); -- 
    minSumDecode_CP_6680_elements(1011) <= minSumDecode_CP_6680_elements(1010);
    -- CP-element group 1012:  merge  place  bypass 
    -- CP-element group 1012: predecessors 
    -- CP-element group 1012: 	1008 
    -- CP-element group 1012: 	1011 
    -- CP-element group 1012: successors 
    -- CP-element group 1012: 	1013 
    -- CP-element group 1012:  members (1) 
      -- CP-element group 1012: 	 branch_block_stmt_1353/merge_stmt_1960_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1012) <= OrReduce(minSumDecode_CP_6680_elements(1008) & minSumDecode_CP_6680_elements(1011));
    -- CP-element group 1013:  transition  bypass 
    -- CP-element group 1013: predecessors 
    -- CP-element group 1013: 	1012 
    -- CP-element group 1013: successors 
    -- CP-element group 1013: 	1014 
    -- CP-element group 1013:  members (1) 
      -- CP-element group 1013: 	 branch_block_stmt_1353/merge_stmt_1960_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1013) <= minSumDecode_CP_6680_elements(1012);
    -- CP-element group 1014:  transition  input  no-bypass 
    -- CP-element group 1014: predecessors 
    -- CP-element group 1014: 	1013 
    -- CP-element group 1014: successors 
    -- CP-element group 1014: 	46 
    -- CP-element group 1014:  members (2) 
      -- CP-element group 1014: 	 branch_block_stmt_1353/merge_stmt_1960_PhiAck/$exit
      -- CP-element group 1014: 	 branch_block_stmt_1353/merge_stmt_1960_PhiAck/phi_stmt_1961_ack
      -- 
    phi_stmt_1961_ack_12647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1014_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1961_ack_0, ack => minSumDecode_CP_6680_elements(1014)); -- 
    -- CP-element group 1015:  transition  bypass 
    -- CP-element group 1015: predecessors 
    -- CP-element group 1015: 	514 
    -- CP-element group 1015: successors 
    -- CP-element group 1015: 	1016 
    -- CP-element group 1015:  members (2) 
      -- CP-element group 1015: 	 branch_block_stmt_1353/bb_24_update_aPosteriorix_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 1015: 	 branch_block_stmt_1353/bb_24_update_aPosteriorix_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1015) <= minSumDecode_CP_6680_elements(514);
    -- CP-element group 1016:  place  bypass 
    -- CP-element group 1016: predecessors 
    -- CP-element group 1016: 	1015 
    -- CP-element group 1016: successors 
    -- CP-element group 1016: 	1017 
    -- CP-element group 1016:  members (1) 
      -- CP-element group 1016: 	 branch_block_stmt_1353/merge_stmt_2038_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1016) <= minSumDecode_CP_6680_elements(1015);
    -- CP-element group 1017:  transition  bypass 
    -- CP-element group 1017: predecessors 
    -- CP-element group 1017: 	1016 
    -- CP-element group 1017: successors 
    -- CP-element group 1017: 	48 
    -- CP-element group 1017:  members (3) 
      -- CP-element group 1017: 	 branch_block_stmt_1353/merge_stmt_2038_PhiAck/$entry
      -- CP-element group 1017: 	 branch_block_stmt_1353/merge_stmt_2038_PhiAck/$exit
      -- CP-element group 1017: 	 branch_block_stmt_1353/merge_stmt_2038_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1017) <= minSumDecode_CP_6680_elements(1016);
    -- CP-element group 1018:  transition  bypass 
    -- CP-element group 1018: predecessors 
    -- CP-element group 1018: 	461 
    -- CP-element group 1018: successors 
    -- CP-element group 1018: 	1020 
    -- CP-element group 1018:  members (2) 
      -- CP-element group 1018: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_update_aPosteriorix_xexit_PhiReq/$entry
      -- CP-element group 1018: 	 branch_block_stmt_1353/initializeExtrinsicInfox_xexit_update_aPosteriorix_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1018) <= minSumDecode_CP_6680_elements(461);
    -- CP-element group 1019:  transition  bypass 
    -- CP-element group 1019: predecessors 
    -- CP-element group 1019: 	48 
    -- CP-element group 1019: successors 
    -- CP-element group 1019: 	1020 
    -- CP-element group 1019:  members (2) 
      -- CP-element group 1019: 	 branch_block_stmt_1353/update_aPosteriorix_xexitx_xloopexit_update_aPosteriorix_xexit_PhiReq/$entry
      -- CP-element group 1019: 	 branch_block_stmt_1353/update_aPosteriorix_xexitx_xloopexit_update_aPosteriorix_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1019) <= minSumDecode_CP_6680_elements(48);
    -- CP-element group 1020:  merge  place  bypass 
    -- CP-element group 1020: predecessors 
    -- CP-element group 1020: 	1018 
    -- CP-element group 1020: 	1019 
    -- CP-element group 1020: successors 
    -- CP-element group 1020: 	1021 
    -- CP-element group 1020:  members (1) 
      -- CP-element group 1020: 	 branch_block_stmt_1353/merge_stmt_2040_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1020) <= OrReduce(minSumDecode_CP_6680_elements(1018) & minSumDecode_CP_6680_elements(1019));
    -- CP-element group 1021:  transition  bypass 
    -- CP-element group 1021: predecessors 
    -- CP-element group 1021: 	1020 
    -- CP-element group 1021: successors 
    -- CP-element group 1021: 	49 
    -- CP-element group 1021:  members (3) 
      -- CP-element group 1021: 	 branch_block_stmt_1353/merge_stmt_2040_PhiAck/$entry
      -- CP-element group 1021: 	 branch_block_stmt_1353/merge_stmt_2040_PhiAck/$exit
      -- CP-element group 1021: 	 branch_block_stmt_1353/merge_stmt_2040_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1021) <= minSumDecode_CP_6680_elements(1020);
    -- CP-element group 1022:  fork  transition  output  bypass 
    -- CP-element group 1022: predecessors 
    -- CP-element group 1022: 	531 
    -- CP-element group 1022: successors 
    -- CP-element group 1022: 	1023 
    -- CP-element group 1022: 	1024 
    -- CP-element group 1022:  members (9) 
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/rr
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/$entry
      -- CP-element group 1022: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/cr
      -- 
    rr_12693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1022), ack => type_cast_2064_inst_req_0); -- 
    cr_12698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1022), ack => type_cast_2064_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1022) <= minSumDecode_CP_6680_elements(531);
    -- CP-element group 1023:  transition  input  no-bypass 
    -- CP-element group 1023: predecessors 
    -- CP-element group 1023: 	1022 
    -- CP-element group 1023: successors 
    -- CP-element group 1023: 	1025 
    -- CP-element group 1023:  members (2) 
      -- CP-element group 1023: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/$exit
      -- CP-element group 1023: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Sample/ra
      -- 
    ra_12694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1023_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_0, ack => minSumDecode_CP_6680_elements(1023)); -- 
    -- CP-element group 1024:  transition  input  no-bypass 
    -- CP-element group 1024: predecessors 
    -- CP-element group 1024: 	1022 
    -- CP-element group 1024: successors 
    -- CP-element group 1024: 	1025 
    -- CP-element group 1024:  members (2) 
      -- CP-element group 1024: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/$exit
      -- CP-element group 1024: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/Update/ca
      -- 
    ca_12699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1024_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_1, ack => minSumDecode_CP_6680_elements(1024)); -- 
    -- CP-element group 1025:  join  transition  output  bypass 
    -- CP-element group 1025: predecessors 
    -- CP-element group 1025: 	1023 
    -- CP-element group 1025: 	1024 
    -- CP-element group 1025: successors 
    -- CP-element group 1025: 	1026 
    -- CP-element group 1025:  members (6) 
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/$exit
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/$exit
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$exit
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/$exit
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2064/SplitProtocol/$exit
      -- CP-element group 1025: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_checkIsdecodedx_xexitx_xthreadx_xthread_PhiReq/phi_stmt_2061/phi_stmt_2061_req
      -- 
    phi_stmt_2061_req_12700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2061_req_12700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1025), ack => phi_stmt_2061_req_0); -- 
    minSumDecode_cp_element_group_1025: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1025"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1023) & minSumDecode_CP_6680_elements(1024);
      gj_minSumDecode_cp_element_group_1025 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1025), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1026:  place  bypass 
    -- CP-element group 1026: predecessors 
    -- CP-element group 1026: 	1025 
    -- CP-element group 1026: successors 
    -- CP-element group 1026: 	1027 
    -- CP-element group 1026:  members (1) 
      -- CP-element group 1026: 	 branch_block_stmt_1353/merge_stmt_2060_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1026) <= minSumDecode_CP_6680_elements(1025);
    -- CP-element group 1027:  transition  bypass 
    -- CP-element group 1027: predecessors 
    -- CP-element group 1027: 	1026 
    -- CP-element group 1027: successors 
    -- CP-element group 1027: 	1028 
    -- CP-element group 1027:  members (1) 
      -- CP-element group 1027: 	 branch_block_stmt_1353/merge_stmt_2060_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1027) <= minSumDecode_CP_6680_elements(1026);
    -- CP-element group 1028:  transition  input  no-bypass 
    -- CP-element group 1028: predecessors 
    -- CP-element group 1028: 	1027 
    -- CP-element group 1028: successors 
    -- CP-element group 1028: 	51 
    -- CP-element group 1028:  members (2) 
      -- CP-element group 1028: 	 branch_block_stmt_1353/merge_stmt_2060_PhiAck/$exit
      -- CP-element group 1028: 	 branch_block_stmt_1353/merge_stmt_2060_PhiAck/phi_stmt_2061_ack
      -- 
    phi_stmt_2061_ack_12705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1028_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2061_ack_0, ack => minSumDecode_CP_6680_elements(1028)); -- 
    -- CP-element group 1029:  transition  bypass 
    -- CP-element group 1029: predecessors 
    -- CP-element group 1029: 	532 
    -- CP-element group 1029: successors 
    -- CP-element group 1029: 	1030 
    -- CP-element group 1029:  members (2) 
      -- CP-element group 1029: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_bbx_xnphx_xi43_PhiReq/$entry
      -- CP-element group 1029: 	 branch_block_stmt_1353/update_aPosteriorix_xexit_bbx_xnphx_xi43_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1029) <= minSumDecode_CP_6680_elements(532);
    -- CP-element group 1030:  place  bypass 
    -- CP-element group 1030: predecessors 
    -- CP-element group 1030: 	1029 
    -- CP-element group 1030: successors 
    -- CP-element group 1030: 	1031 
    -- CP-element group 1030:  members (1) 
      -- CP-element group 1030: 	 branch_block_stmt_1353/merge_stmt_2070_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1030) <= minSumDecode_CP_6680_elements(1029);
    -- CP-element group 1031:  transition  bypass 
    -- CP-element group 1031: predecessors 
    -- CP-element group 1031: 	1030 
    -- CP-element group 1031: successors 
    -- CP-element group 1031: 	53 
    -- CP-element group 1031:  members (3) 
      -- CP-element group 1031: 	 branch_block_stmt_1353/merge_stmt_2070_PhiAck/$entry
      -- CP-element group 1031: 	 branch_block_stmt_1353/merge_stmt_2070_PhiAck/$exit
      -- CP-element group 1031: 	 branch_block_stmt_1353/merge_stmt_2070_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1031) <= minSumDecode_CP_6680_elements(1030);
    -- CP-element group 1032:  fork  transition  output  bypass 
    -- CP-element group 1032: predecessors 
    -- CP-element group 1032: 	639 
    -- CP-element group 1032: successors 
    -- CP-element group 1032: 	1033 
    -- CP-element group 1032: 	1034 
    -- CP-element group 1032: 	1036 
    -- CP-element group 1032: 	1037 
    -- CP-element group 1032:  members (17) 
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Sample/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Sample/rr
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Update/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Update/cr
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Sample/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Sample/rr
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Update/$entry
      -- CP-element group 1032: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Update/cr
      -- 
    rr_12732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1032), ack => type_cast_2115_inst_req_0); -- 
    cr_12737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1032), ack => type_cast_2115_inst_req_1); -- 
    rr_12755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1032), ack => type_cast_2108_inst_req_0); -- 
    cr_12760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1032), ack => type_cast_2108_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1032) <= minSumDecode_CP_6680_elements(639);
    -- CP-element group 1033:  transition  input  no-bypass 
    -- CP-element group 1033: predecessors 
    -- CP-element group 1033: 	1032 
    -- CP-element group 1033: successors 
    -- CP-element group 1033: 	1035 
    -- CP-element group 1033:  members (2) 
      -- CP-element group 1033: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Sample/$exit
      -- CP-element group 1033: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Sample/ra
      -- 
    ra_12733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1033_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2115_inst_ack_0, ack => minSumDecode_CP_6680_elements(1033)); -- 
    -- CP-element group 1034:  transition  input  no-bypass 
    -- CP-element group 1034: predecessors 
    -- CP-element group 1034: 	1032 
    -- CP-element group 1034: successors 
    -- CP-element group 1034: 	1035 
    -- CP-element group 1034:  members (2) 
      -- CP-element group 1034: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Update/$exit
      -- CP-element group 1034: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/Update/ca
      -- 
    ca_12738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1034_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2115_inst_ack_1, ack => minSumDecode_CP_6680_elements(1034)); -- 
    -- CP-element group 1035:  join  transition  output  bypass 
    -- CP-element group 1035: predecessors 
    -- CP-element group 1035: 	1033 
    -- CP-element group 1035: 	1034 
    -- CP-element group 1035: successors 
    -- CP-element group 1035: 	1039 
    -- CP-element group 1035:  members (5) 
      -- CP-element group 1035: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/$exit
      -- CP-element group 1035: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/$exit
      -- CP-element group 1035: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/$exit
      -- CP-element group 1035: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2115/SplitProtocol/$exit
      -- CP-element group 1035: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_req
      -- 
    phi_stmt_2109_req_12739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2109_req_12739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1035), ack => phi_stmt_2109_req_1); -- 
    minSumDecode_cp_element_group_1035: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1035"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1033) & minSumDecode_CP_6680_elements(1034);
      gj_minSumDecode_cp_element_group_1035 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1035), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1036:  transition  input  no-bypass 
    -- CP-element group 1036: predecessors 
    -- CP-element group 1036: 	1032 
    -- CP-element group 1036: successors 
    -- CP-element group 1036: 	1038 
    -- CP-element group 1036:  members (2) 
      -- CP-element group 1036: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Sample/$exit
      -- CP-element group 1036: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Sample/ra
      -- 
    ra_12756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1036_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2108_inst_ack_0, ack => minSumDecode_CP_6680_elements(1036)); -- 
    -- CP-element group 1037:  transition  input  no-bypass 
    -- CP-element group 1037: predecessors 
    -- CP-element group 1037: 	1032 
    -- CP-element group 1037: successors 
    -- CP-element group 1037: 	1038 
    -- CP-element group 1037:  members (2) 
      -- CP-element group 1037: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Update/$exit
      -- CP-element group 1037: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/Update/ca
      -- 
    ca_12761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1037_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2108_inst_ack_1, ack => minSumDecode_CP_6680_elements(1037)); -- 
    -- CP-element group 1038:  join  transition  output  bypass 
    -- CP-element group 1038: predecessors 
    -- CP-element group 1038: 	1036 
    -- CP-element group 1038: 	1037 
    -- CP-element group 1038: successors 
    -- CP-element group 1038: 	1039 
    -- CP-element group 1038:  members (5) 
      -- CP-element group 1038: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/$exit
      -- CP-element group 1038: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/$exit
      -- CP-element group 1038: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/$exit
      -- CP-element group 1038: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2108/SplitProtocol/$exit
      -- CP-element group 1038: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_req
      -- 
    phi_stmt_2102_req_12762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2102_req_12762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1038), ack => phi_stmt_2102_req_1); -- 
    minSumDecode_cp_element_group_1038: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1038"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1036) & minSumDecode_CP_6680_elements(1037);
      gj_minSumDecode_cp_element_group_1038 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1038), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1039:  join  transition  bypass 
    -- CP-element group 1039: predecessors 
    -- CP-element group 1039: 	1035 
    -- CP-element group 1039: 	1038 
    -- CP-element group 1039: successors 
    -- CP-element group 1039: 	1046 
    -- CP-element group 1039:  members (1) 
      -- CP-element group 1039: 	 branch_block_stmt_1353/bb_37_bb_29_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1039: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1039"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1035) & minSumDecode_CP_6680_elements(1038);
      gj_minSumDecode_cp_element_group_1039 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1039), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1040:  fork  transition  bypass 
    -- CP-element group 1040: predecessors 
    -- CP-element group 1040: 	54 
    -- CP-element group 1040: successors 
    -- CP-element group 1040: 	1041 
    -- CP-element group 1040: 	1043 
    -- CP-element group 1040:  members (5) 
      -- CP-element group 1040: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/$entry
      -- CP-element group 1040: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/$entry
      -- CP-element group 1040: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/$entry
      -- CP-element group 1040: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/$entry
      -- CP-element group 1040: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1040) <= minSumDecode_CP_6680_elements(54);
    -- CP-element group 1041:  transition  bypass 
    -- CP-element group 1041: predecessors 
    -- CP-element group 1041: 	1040 
    -- CP-element group 1041: successors 
    -- CP-element group 1041: 	1042 
    -- CP-element group 1041:  members (1) 
      -- CP-element group 1041: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/type_cast_2113_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1041) is a control-delay.
    cp_element_1041_delay: control_delay_element  generic map(name => " 1041_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1040), ack => minSumDecode_CP_6680_elements(1041), clk => clk, reset =>reset);
    -- CP-element group 1042:  transition  output  bypass 
    -- CP-element group 1042: predecessors 
    -- CP-element group 1042: 	1041 
    -- CP-element group 1042: successors 
    -- CP-element group 1042: 	1045 
    -- CP-element group 1042:  members (3) 
      -- CP-element group 1042: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/$exit
      -- CP-element group 1042: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_sources/$exit
      -- CP-element group 1042: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2109/phi_stmt_2109_req
      -- 
    phi_stmt_2109_req_12773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2109_req_12773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1042), ack => phi_stmt_2109_req_0); -- 
    minSumDecode_CP_6680_elements(1042) <= minSumDecode_CP_6680_elements(1041);
    -- CP-element group 1043:  transition  bypass 
    -- CP-element group 1043: predecessors 
    -- CP-element group 1043: 	1040 
    -- CP-element group 1043: successors 
    -- CP-element group 1043: 	1044 
    -- CP-element group 1043:  members (1) 
      -- CP-element group 1043: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/type_cast_2106_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1043) is a control-delay.
    cp_element_1043_delay: control_delay_element  generic map(name => " 1043_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1040), ack => minSumDecode_CP_6680_elements(1043), clk => clk, reset =>reset);
    -- CP-element group 1044:  transition  output  bypass 
    -- CP-element group 1044: predecessors 
    -- CP-element group 1044: 	1043 
    -- CP-element group 1044: successors 
    -- CP-element group 1044: 	1045 
    -- CP-element group 1044:  members (3) 
      -- CP-element group 1044: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/$exit
      -- CP-element group 1044: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_sources/$exit
      -- CP-element group 1044: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/phi_stmt_2102/phi_stmt_2102_req
      -- 
    phi_stmt_2102_req_12781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2102_req_12781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1044), ack => phi_stmt_2102_req_0); -- 
    minSumDecode_CP_6680_elements(1044) <= minSumDecode_CP_6680_elements(1043);
    -- CP-element group 1045:  join  transition  no-bypass 
    -- CP-element group 1045: predecessors 
    -- CP-element group 1045: 	1042 
    -- CP-element group 1045: 	1044 
    -- CP-element group 1045: successors 
    -- CP-element group 1045: 	1046 
    -- CP-element group 1045:  members (1) 
      -- CP-element group 1045: 	 branch_block_stmt_1353/bbx_xnphx_xi43_bb_29_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1045: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1045"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1042) & minSumDecode_CP_6680_elements(1044);
      gj_minSumDecode_cp_element_group_1045 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1045), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1046:  merge  place  bypass 
    -- CP-element group 1046: predecessors 
    -- CP-element group 1046: 	1039 
    -- CP-element group 1046: 	1045 
    -- CP-element group 1046: successors 
    -- CP-element group 1046: 	1047 
    -- CP-element group 1046:  members (1) 
      -- CP-element group 1046: 	 branch_block_stmt_1353/merge_stmt_2101_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1046) <= OrReduce(minSumDecode_CP_6680_elements(1039) & minSumDecode_CP_6680_elements(1045));
    -- CP-element group 1047:  fork  transition  bypass 
    -- CP-element group 1047: predecessors 
    -- CP-element group 1047: 	1046 
    -- CP-element group 1047: successors 
    -- CP-element group 1047: 	1048 
    -- CP-element group 1047: 	1049 
    -- CP-element group 1047:  members (1) 
      -- CP-element group 1047: 	 branch_block_stmt_1353/merge_stmt_2101_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1047) <= minSumDecode_CP_6680_elements(1046);
    -- CP-element group 1048:  transition  input  no-bypass 
    -- CP-element group 1048: predecessors 
    -- CP-element group 1048: 	1047 
    -- CP-element group 1048: successors 
    -- CP-element group 1048: 	1050 
    -- CP-element group 1048:  members (1) 
      -- CP-element group 1048: 	 branch_block_stmt_1353/merge_stmt_2101_PhiAck/phi_stmt_2102_ack
      -- 
    phi_stmt_2102_ack_12786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1048_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2102_ack_0, ack => minSumDecode_CP_6680_elements(1048)); -- 
    -- CP-element group 1049:  transition  input  no-bypass 
    -- CP-element group 1049: predecessors 
    -- CP-element group 1049: 	1047 
    -- CP-element group 1049: successors 
    -- CP-element group 1049: 	1050 
    -- CP-element group 1049:  members (1) 
      -- CP-element group 1049: 	 branch_block_stmt_1353/merge_stmt_2101_PhiAck/phi_stmt_2109_ack
      -- 
    phi_stmt_2109_ack_12787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1049_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2109_ack_0, ack => minSumDecode_CP_6680_elements(1049)); -- 
    -- CP-element group 1050:  join  transition  bypass 
    -- CP-element group 1050: predecessors 
    -- CP-element group 1050: 	1048 
    -- CP-element group 1050: 	1049 
    -- CP-element group 1050: successors 
    -- CP-element group 1050: 	55 
    -- CP-element group 1050:  members (1) 
      -- CP-element group 1050: 	 branch_block_stmt_1353/merge_stmt_2101_PhiAck/$exit
      -- 
    minSumDecode_cp_element_group_1050: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1050"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1048) & minSumDecode_CP_6680_elements(1049);
      gj_minSumDecode_cp_element_group_1050 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1050), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1051:  transition  bypass 
    -- CP-element group 1051: predecessors 
    -- CP-element group 1051: 	568 
    -- CP-element group 1051: successors 
    -- CP-element group 1051: 	1052 
    -- CP-element group 1051:  members (2) 
      -- CP-element group 1051: 	 branch_block_stmt_1353/bb_29_bb_30_PhiReq/$entry
      -- CP-element group 1051: 	 branch_block_stmt_1353/bb_29_bb_30_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1051) <= minSumDecode_CP_6680_elements(568);
    -- CP-element group 1052:  place  bypass 
    -- CP-element group 1052: predecessors 
    -- CP-element group 1052: 	1051 
    -- CP-element group 1052: successors 
    -- CP-element group 1052: 	1053 
    -- CP-element group 1052:  members (1) 
      -- CP-element group 1052: 	 branch_block_stmt_1353/merge_stmt_2147_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1052) <= minSumDecode_CP_6680_elements(1051);
    -- CP-element group 1053:  transition  bypass 
    -- CP-element group 1053: predecessors 
    -- CP-element group 1053: 	1052 
    -- CP-element group 1053: successors 
    -- CP-element group 1053: 	57 
    -- CP-element group 1053:  members (3) 
      -- CP-element group 1053: 	 branch_block_stmt_1353/merge_stmt_2147_PhiAck/$entry
      -- CP-element group 1053: 	 branch_block_stmt_1353/merge_stmt_2147_PhiAck/$exit
      -- CP-element group 1053: 	 branch_block_stmt_1353/merge_stmt_2147_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1053) <= minSumDecode_CP_6680_elements(1052);
    -- CP-element group 1054:  transition  bypass 
    -- CP-element group 1054: predecessors 
    -- CP-element group 1054: 	584 
    -- CP-element group 1054: successors 
    -- CP-element group 1054: 	1055 
    -- CP-element group 1054:  members (2) 
      -- CP-element group 1054: 	 branch_block_stmt_1353/bb_30_bb_31_PhiReq/$entry
      -- CP-element group 1054: 	 branch_block_stmt_1353/bb_30_bb_31_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1054) <= minSumDecode_CP_6680_elements(584);
    -- CP-element group 1055:  place  bypass 
    -- CP-element group 1055: predecessors 
    -- CP-element group 1055: 	1054 
    -- CP-element group 1055: successors 
    -- CP-element group 1055: 	1056 
    -- CP-element group 1055:  members (1) 
      -- CP-element group 1055: 	 branch_block_stmt_1353/merge_stmt_2168_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1055) <= minSumDecode_CP_6680_elements(1054);
    -- CP-element group 1056:  transition  bypass 
    -- CP-element group 1056: predecessors 
    -- CP-element group 1056: 	1055 
    -- CP-element group 1056: successors 
    -- CP-element group 1056: 	59 
    -- CP-element group 1056:  members (3) 
      -- CP-element group 1056: 	 branch_block_stmt_1353/merge_stmt_2168_PhiAck/$entry
      -- CP-element group 1056: 	 branch_block_stmt_1353/merge_stmt_2168_PhiAck/$exit
      -- CP-element group 1056: 	 branch_block_stmt_1353/merge_stmt_2168_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1056) <= minSumDecode_CP_6680_elements(1055);
    -- CP-element group 1057:  fork  transition  output  bypass 
    -- CP-element group 1057: predecessors 
    -- CP-element group 1057: 	585 
    -- CP-element group 1057: successors 
    -- CP-element group 1057: 	1058 
    -- CP-element group 1057: 	1059 
    -- CP-element group 1057:  members (9) 
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/rr
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/$entry
      -- CP-element group 1057: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/cr
      -- 
    rr_12830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1057), ack => type_cast_2181_inst_req_0); -- 
    cr_12835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1057), ack => type_cast_2181_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1057) <= minSumDecode_CP_6680_elements(585);
    -- CP-element group 1058:  transition  input  no-bypass 
    -- CP-element group 1058: predecessors 
    -- CP-element group 1058: 	1057 
    -- CP-element group 1058: successors 
    -- CP-element group 1058: 	1060 
    -- CP-element group 1058:  members (2) 
      -- CP-element group 1058: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/$exit
      -- CP-element group 1058: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Sample/ra
      -- 
    ra_12831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1058_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_0, ack => minSumDecode_CP_6680_elements(1058)); -- 
    -- CP-element group 1059:  transition  input  no-bypass 
    -- CP-element group 1059: predecessors 
    -- CP-element group 1059: 	1057 
    -- CP-element group 1059: successors 
    -- CP-element group 1059: 	1060 
    -- CP-element group 1059:  members (2) 
      -- CP-element group 1059: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/$exit
      -- CP-element group 1059: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/Update/ca
      -- 
    ca_12836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1059_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_1, ack => minSumDecode_CP_6680_elements(1059)); -- 
    -- CP-element group 1060:  join  transition  output  bypass 
    -- CP-element group 1060: predecessors 
    -- CP-element group 1060: 	1058 
    -- CP-element group 1060: 	1059 
    -- CP-element group 1060: successors 
    -- CP-element group 1060: 	1064 
    -- CP-element group 1060:  members (6) 
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/$exit
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/$exit
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/$exit
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2181/SplitProtocol/$exit
      -- CP-element group 1060: 	 branch_block_stmt_1353/bb_30_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- 
    phi_stmt_2175_req_12837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_12837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1060), ack => phi_stmt_2175_req_1); -- 
    minSumDecode_cp_element_group_1060: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1060"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1058) & minSumDecode_CP_6680_elements(1059);
      gj_minSumDecode_cp_element_group_1060 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1060), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1061:  transition  bypass 
    -- CP-element group 1061: predecessors 
    -- CP-element group 1061: 	60 
    -- CP-element group 1061: successors 
    -- CP-element group 1061: 	1062 
    -- CP-element group 1061:  members (3) 
      -- CP-element group 1061: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/$entry
      -- CP-element group 1061: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/$entry
      -- CP-element group 1061: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1061) <= minSumDecode_CP_6680_elements(60);
    -- CP-element group 1062:  transition  bypass 
    -- CP-element group 1062: predecessors 
    -- CP-element group 1062: 	1061 
    -- CP-element group 1062: successors 
    -- CP-element group 1062: 	1063 
    -- CP-element group 1062:  members (1) 
      -- CP-element group 1062: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/type_cast_2179_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1062) is a control-delay.
    cp_element_1062_delay: control_delay_element  generic map(name => " 1062_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1061), ack => minSumDecode_CP_6680_elements(1062), clk => clk, reset =>reset);
    -- CP-element group 1063:  transition  output  bypass 
    -- CP-element group 1063: predecessors 
    -- CP-element group 1063: 	1062 
    -- CP-element group 1063: successors 
    -- CP-element group 1063: 	1064 
    -- CP-element group 1063:  members (4) 
      -- CP-element group 1063: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/$exit
      -- CP-element group 1063: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/$exit
      -- CP-element group 1063: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_sources/$exit
      -- CP-element group 1063: 	 branch_block_stmt_1353/bb_31_bb_32_PhiReq/phi_stmt_2175/phi_stmt_2175_req
      -- 
    phi_stmt_2175_req_12848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2175_req_12848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1063), ack => phi_stmt_2175_req_0); -- 
    minSumDecode_CP_6680_elements(1063) <= minSumDecode_CP_6680_elements(1062);
    -- CP-element group 1064:  merge  place  bypass 
    -- CP-element group 1064: predecessors 
    -- CP-element group 1064: 	1060 
    -- CP-element group 1064: 	1063 
    -- CP-element group 1064: successors 
    -- CP-element group 1064: 	1065 
    -- CP-element group 1064:  members (1) 
      -- CP-element group 1064: 	 branch_block_stmt_1353/merge_stmt_2174_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1064) <= OrReduce(minSumDecode_CP_6680_elements(1060) & minSumDecode_CP_6680_elements(1063));
    -- CP-element group 1065:  transition  bypass 
    -- CP-element group 1065: predecessors 
    -- CP-element group 1065: 	1064 
    -- CP-element group 1065: successors 
    -- CP-element group 1065: 	1066 
    -- CP-element group 1065:  members (1) 
      -- CP-element group 1065: 	 branch_block_stmt_1353/merge_stmt_2174_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1065) <= minSumDecode_CP_6680_elements(1064);
    -- CP-element group 1066:  transition  input  no-bypass 
    -- CP-element group 1066: predecessors 
    -- CP-element group 1066: 	1065 
    -- CP-element group 1066: successors 
    -- CP-element group 1066: 	61 
    -- CP-element group 1066:  members (2) 
      -- CP-element group 1066: 	 branch_block_stmt_1353/merge_stmt_2174_PhiAck/$exit
      -- CP-element group 1066: 	 branch_block_stmt_1353/merge_stmt_2174_PhiAck/phi_stmt_2175_ack
      -- 
    phi_stmt_2175_ack_12853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1066_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2175_ack_0, ack => minSumDecode_CP_6680_elements(1066)); -- 
    -- CP-element group 1067:  transition  bypass 
    -- CP-element group 1067: predecessors 
    -- CP-element group 1067: 	569 
    -- CP-element group 1067: successors 
    -- CP-element group 1067: 	1068 
    -- CP-element group 1067:  members (2) 
      -- CP-element group 1067: 	 branch_block_stmt_1353/bb_29_bb_33_PhiReq/$entry
      -- CP-element group 1067: 	 branch_block_stmt_1353/bb_29_bb_33_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1067) <= minSumDecode_CP_6680_elements(569);
    -- CP-element group 1068:  place  bypass 
    -- CP-element group 1068: predecessors 
    -- CP-element group 1068: 	1067 
    -- CP-element group 1068: successors 
    -- CP-element group 1068: 	1069 
    -- CP-element group 1068:  members (1) 
      -- CP-element group 1068: 	 branch_block_stmt_1353/merge_stmt_2189_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1068) <= minSumDecode_CP_6680_elements(1067);
    -- CP-element group 1069:  transition  bypass 
    -- CP-element group 1069: predecessors 
    -- CP-element group 1069: 	1068 
    -- CP-element group 1069: successors 
    -- CP-element group 1069: 	63 
    -- CP-element group 1069:  members (3) 
      -- CP-element group 1069: 	 branch_block_stmt_1353/merge_stmt_2189_PhiAck/$entry
      -- CP-element group 1069: 	 branch_block_stmt_1353/merge_stmt_2189_PhiAck/$exit
      -- CP-element group 1069: 	 branch_block_stmt_1353/merge_stmt_2189_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1069) <= minSumDecode_CP_6680_elements(1068);
    -- CP-element group 1070:  transition  bypass 
    -- CP-element group 1070: predecessors 
    -- CP-element group 1070: 	602 
    -- CP-element group 1070: successors 
    -- CP-element group 1070: 	1071 
    -- CP-element group 1070:  members (2) 
      -- CP-element group 1070: 	 branch_block_stmt_1353/bb_33_bb_34_PhiReq/$entry
      -- CP-element group 1070: 	 branch_block_stmt_1353/bb_33_bb_34_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1070) <= minSumDecode_CP_6680_elements(602);
    -- CP-element group 1071:  place  bypass 
    -- CP-element group 1071: predecessors 
    -- CP-element group 1071: 	1070 
    -- CP-element group 1071: successors 
    -- CP-element group 1071: 	1072 
    -- CP-element group 1071:  members (1) 
      -- CP-element group 1071: 	 branch_block_stmt_1353/merge_stmt_2202_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1071) <= minSumDecode_CP_6680_elements(1070);
    -- CP-element group 1072:  transition  bypass 
    -- CP-element group 1072: predecessors 
    -- CP-element group 1072: 	1071 
    -- CP-element group 1072: successors 
    -- CP-element group 1072: 	65 
    -- CP-element group 1072:  members (3) 
      -- CP-element group 1072: 	 branch_block_stmt_1353/merge_stmt_2202_PhiAck/$entry
      -- CP-element group 1072: 	 branch_block_stmt_1353/merge_stmt_2202_PhiAck/$exit
      -- CP-element group 1072: 	 branch_block_stmt_1353/merge_stmt_2202_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1072) <= minSumDecode_CP_6680_elements(1071);
    -- CP-element group 1073:  transition  bypass 
    -- CP-element group 1073: predecessors 
    -- CP-element group 1073: 	618 
    -- CP-element group 1073: successors 
    -- CP-element group 1073: 	1074 
    -- CP-element group 1073:  members (2) 
      -- CP-element group 1073: 	 branch_block_stmt_1353/bb_34_bb_35_PhiReq/$entry
      -- CP-element group 1073: 	 branch_block_stmt_1353/bb_34_bb_35_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1073) <= minSumDecode_CP_6680_elements(618);
    -- CP-element group 1074:  place  bypass 
    -- CP-element group 1074: predecessors 
    -- CP-element group 1074: 	1073 
    -- CP-element group 1074: successors 
    -- CP-element group 1074: 	1075 
    -- CP-element group 1074:  members (1) 
      -- CP-element group 1074: 	 branch_block_stmt_1353/merge_stmt_2223_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1074) <= minSumDecode_CP_6680_elements(1073);
    -- CP-element group 1075:  transition  bypass 
    -- CP-element group 1075: predecessors 
    -- CP-element group 1075: 	1074 
    -- CP-element group 1075: successors 
    -- CP-element group 1075: 	67 
    -- CP-element group 1075:  members (3) 
      -- CP-element group 1075: 	 branch_block_stmt_1353/merge_stmt_2223_PhiAck/$entry
      -- CP-element group 1075: 	 branch_block_stmt_1353/merge_stmt_2223_PhiAck/$exit
      -- CP-element group 1075: 	 branch_block_stmt_1353/merge_stmt_2223_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1075) <= minSumDecode_CP_6680_elements(1074);
    -- CP-element group 1076:  fork  transition  output  bypass 
    -- CP-element group 1076: predecessors 
    -- CP-element group 1076: 	619 
    -- CP-element group 1076: successors 
    -- CP-element group 1076: 	1077 
    -- CP-element group 1076: 	1078 
    -- CP-element group 1076:  members (9) 
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Sample/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Sample/rr
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Update/$entry
      -- CP-element group 1076: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Update/cr
      -- 
    rr_12904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1076), ack => type_cast_2236_inst_req_0); -- 
    cr_12909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1076), ack => type_cast_2236_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1076) <= minSumDecode_CP_6680_elements(619);
    -- CP-element group 1077:  transition  input  no-bypass 
    -- CP-element group 1077: predecessors 
    -- CP-element group 1077: 	1076 
    -- CP-element group 1077: successors 
    -- CP-element group 1077: 	1079 
    -- CP-element group 1077:  members (2) 
      -- CP-element group 1077: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Sample/$exit
      -- CP-element group 1077: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Sample/ra
      -- 
    ra_12905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1077_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2236_inst_ack_0, ack => minSumDecode_CP_6680_elements(1077)); -- 
    -- CP-element group 1078:  transition  input  no-bypass 
    -- CP-element group 1078: predecessors 
    -- CP-element group 1078: 	1076 
    -- CP-element group 1078: successors 
    -- CP-element group 1078: 	1079 
    -- CP-element group 1078:  members (2) 
      -- CP-element group 1078: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Update/$exit
      -- CP-element group 1078: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/Update/ca
      -- 
    ca_12910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1078_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2236_inst_ack_1, ack => minSumDecode_CP_6680_elements(1078)); -- 
    -- CP-element group 1079:  join  transition  output  bypass 
    -- CP-element group 1079: predecessors 
    -- CP-element group 1079: 	1077 
    -- CP-element group 1079: 	1078 
    -- CP-element group 1079: successors 
    -- CP-element group 1079: 	1083 
    -- CP-element group 1079:  members (6) 
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/$exit
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/$exit
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/$exit
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/$exit
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2236/SplitProtocol/$exit
      -- CP-element group 1079: 	 branch_block_stmt_1353/bb_34_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_req
      -- 
    phi_stmt_2230_req_12911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2230_req_12911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1079), ack => phi_stmt_2230_req_1); -- 
    minSumDecode_cp_element_group_1079: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1079"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1077) & minSumDecode_CP_6680_elements(1078);
      gj_minSumDecode_cp_element_group_1079 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1079), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1080:  transition  bypass 
    -- CP-element group 1080: predecessors 
    -- CP-element group 1080: 	68 
    -- CP-element group 1080: successors 
    -- CP-element group 1080: 	1081 
    -- CP-element group 1080:  members (3) 
      -- CP-element group 1080: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/$entry
      -- CP-element group 1080: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/$entry
      -- CP-element group 1080: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1080) <= minSumDecode_CP_6680_elements(68);
    -- CP-element group 1081:  transition  bypass 
    -- CP-element group 1081: predecessors 
    -- CP-element group 1081: 	1080 
    -- CP-element group 1081: successors 
    -- CP-element group 1081: 	1082 
    -- CP-element group 1081:  members (1) 
      -- CP-element group 1081: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/type_cast_2234_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1081) is a control-delay.
    cp_element_1081_delay: control_delay_element  generic map(name => " 1081_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1080), ack => minSumDecode_CP_6680_elements(1081), clk => clk, reset =>reset);
    -- CP-element group 1082:  transition  output  bypass 
    -- CP-element group 1082: predecessors 
    -- CP-element group 1082: 	1081 
    -- CP-element group 1082: successors 
    -- CP-element group 1082: 	1083 
    -- CP-element group 1082:  members (4) 
      -- CP-element group 1082: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/$exit
      -- CP-element group 1082: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/$exit
      -- CP-element group 1082: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_sources/$exit
      -- CP-element group 1082: 	 branch_block_stmt_1353/bb_35_bb_36_PhiReq/phi_stmt_2230/phi_stmt_2230_req
      -- 
    phi_stmt_2230_req_12922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2230_req_12922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1082), ack => phi_stmt_2230_req_0); -- 
    minSumDecode_CP_6680_elements(1082) <= minSumDecode_CP_6680_elements(1081);
    -- CP-element group 1083:  merge  place  bypass 
    -- CP-element group 1083: predecessors 
    -- CP-element group 1083: 	1079 
    -- CP-element group 1083: 	1082 
    -- CP-element group 1083: successors 
    -- CP-element group 1083: 	1084 
    -- CP-element group 1083:  members (1) 
      -- CP-element group 1083: 	 branch_block_stmt_1353/merge_stmt_2229_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1083) <= OrReduce(minSumDecode_CP_6680_elements(1079) & minSumDecode_CP_6680_elements(1082));
    -- CP-element group 1084:  transition  bypass 
    -- CP-element group 1084: predecessors 
    -- CP-element group 1084: 	1083 
    -- CP-element group 1084: successors 
    -- CP-element group 1084: 	1085 
    -- CP-element group 1084:  members (1) 
      -- CP-element group 1084: 	 branch_block_stmt_1353/merge_stmt_2229_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1084) <= minSumDecode_CP_6680_elements(1083);
    -- CP-element group 1085:  transition  input  no-bypass 
    -- CP-element group 1085: predecessors 
    -- CP-element group 1085: 	1084 
    -- CP-element group 1085: successors 
    -- CP-element group 1085: 	69 
    -- CP-element group 1085:  members (2) 
      -- CP-element group 1085: 	 branch_block_stmt_1353/merge_stmt_2229_PhiAck/phi_stmt_2230_ack
      -- CP-element group 1085: 	 branch_block_stmt_1353/merge_stmt_2229_PhiAck/$exit
      -- 
    phi_stmt_2230_ack_12927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1085_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2230_ack_0, ack => minSumDecode_CP_6680_elements(1085)); -- 
    -- CP-element group 1086:  fork  transition  output  bypass 
    -- CP-element group 1086: predecessors 
    -- CP-element group 1086: 	62 
    -- CP-element group 1086: successors 
    -- CP-element group 1086: 	1087 
    -- CP-element group 1086: 	1088 
    -- CP-element group 1086:  members (9) 
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Update/cr
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Update/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Sample/rr
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Sample/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/$entry
      -- CP-element group 1086: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/$entry
      -- 
    rr_12946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1086), ack => type_cast_2252_inst_req_0); -- 
    cr_12951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1086), ack => type_cast_2252_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1086) <= minSumDecode_CP_6680_elements(62);
    -- CP-element group 1087:  transition  input  no-bypass 
    -- CP-element group 1087: predecessors 
    -- CP-element group 1087: 	1086 
    -- CP-element group 1087: successors 
    -- CP-element group 1087: 	1089 
    -- CP-element group 1087:  members (2) 
      -- CP-element group 1087: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Sample/ra
      -- CP-element group 1087: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Sample/$exit
      -- 
    ra_12947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1087_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_0, ack => minSumDecode_CP_6680_elements(1087)); -- 
    -- CP-element group 1088:  transition  input  no-bypass 
    -- CP-element group 1088: predecessors 
    -- CP-element group 1088: 	1086 
    -- CP-element group 1088: successors 
    -- CP-element group 1088: 	1089 
    -- CP-element group 1088:  members (2) 
      -- CP-element group 1088: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Update/ca
      -- CP-element group 1088: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/Update/$exit
      -- 
    ca_12952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1088_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_1, ack => minSumDecode_CP_6680_elements(1088)); -- 
    -- CP-element group 1089:  join  transition  output  bypass 
    -- CP-element group 1089: predecessors 
    -- CP-element group 1089: 	1087 
    -- CP-element group 1089: 	1088 
    -- CP-element group 1089: successors 
    -- CP-element group 1089: 	1098 
    -- CP-element group 1089:  members (6) 
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_req
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/SplitProtocol/$exit
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2252/$exit
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$exit
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/phi_stmt_2245/$exit
      -- CP-element group 1089: 	 branch_block_stmt_1353/bb_32_bb_37_PhiReq/$exit
      -- 
    phi_stmt_2245_req_12953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2245_req_12953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1089), ack => phi_stmt_2245_req_2); -- 
    minSumDecode_cp_element_group_1089: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1089"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1087) & minSumDecode_CP_6680_elements(1088);
      gj_minSumDecode_cp_element_group_1089 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1089), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1090:  fork  transition  output  bypass 
    -- CP-element group 1090: predecessors 
    -- CP-element group 1090: 	603 
    -- CP-element group 1090: successors 
    -- CP-element group 1090: 	1091 
    -- CP-element group 1090: 	1092 
    -- CP-element group 1090:  members (9) 
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/rr
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/cr
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/$entry
      -- CP-element group 1090: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/$entry
      -- 
    rr_12972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1090), ack => type_cast_2250_inst_req_0); -- 
    cr_12977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1090), ack => type_cast_2250_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1090) <= minSumDecode_CP_6680_elements(603);
    -- CP-element group 1091:  transition  input  no-bypass 
    -- CP-element group 1091: predecessors 
    -- CP-element group 1091: 	1090 
    -- CP-element group 1091: successors 
    -- CP-element group 1091: 	1093 
    -- CP-element group 1091:  members (2) 
      -- CP-element group 1091: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/ra
      -- CP-element group 1091: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/$exit
      -- 
    ra_12973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1091_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_0, ack => minSumDecode_CP_6680_elements(1091)); -- 
    -- CP-element group 1092:  transition  input  no-bypass 
    -- CP-element group 1092: predecessors 
    -- CP-element group 1092: 	1090 
    -- CP-element group 1092: successors 
    -- CP-element group 1092: 	1093 
    -- CP-element group 1092:  members (2) 
      -- CP-element group 1092: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/ca
      -- CP-element group 1092: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/$exit
      -- 
    ca_12978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1092_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_1, ack => minSumDecode_CP_6680_elements(1092)); -- 
    -- CP-element group 1093:  join  transition  output  bypass 
    -- CP-element group 1093: predecessors 
    -- CP-element group 1093: 	1091 
    -- CP-element group 1093: 	1092 
    -- CP-element group 1093: successors 
    -- CP-element group 1093: 	1098 
    -- CP-element group 1093:  members (6) 
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/$exit
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_req
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/$exit
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$exit
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/phi_stmt_2245/$exit
      -- CP-element group 1093: 	 branch_block_stmt_1353/bb_33_bb_37_PhiReq/$exit
      -- 
    phi_stmt_2245_req_12979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2245_req_12979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1093), ack => phi_stmt_2245_req_1); -- 
    minSumDecode_cp_element_group_1093: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1093"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1091) & minSumDecode_CP_6680_elements(1092);
      gj_minSumDecode_cp_element_group_1093 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1093), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1094:  fork  transition  output  bypass 
    -- CP-element group 1094: predecessors 
    -- CP-element group 1094: 	70 
    -- CP-element group 1094: successors 
    -- CP-element group 1094: 	1095 
    -- CP-element group 1094: 	1096 
    -- CP-element group 1094:  members (9) 
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/cr
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/rr
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$entry
      -- CP-element group 1094: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/$entry
      -- 
    rr_12998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1094), ack => type_cast_2248_inst_req_0); -- 
    cr_13003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1094), ack => type_cast_2248_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1094) <= minSumDecode_CP_6680_elements(70);
    -- CP-element group 1095:  transition  input  no-bypass 
    -- CP-element group 1095: predecessors 
    -- CP-element group 1095: 	1094 
    -- CP-element group 1095: successors 
    -- CP-element group 1095: 	1097 
    -- CP-element group 1095:  members (2) 
      -- CP-element group 1095: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/ra
      -- CP-element group 1095: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/$exit
      -- 
    ra_12999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1095_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_0, ack => minSumDecode_CP_6680_elements(1095)); -- 
    -- CP-element group 1096:  transition  input  no-bypass 
    -- CP-element group 1096: predecessors 
    -- CP-element group 1096: 	1094 
    -- CP-element group 1096: successors 
    -- CP-element group 1096: 	1097 
    -- CP-element group 1096:  members (2) 
      -- CP-element group 1096: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/ca
      -- CP-element group 1096: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/$exit
      -- 
    ca_13004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1096_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_1, ack => minSumDecode_CP_6680_elements(1096)); -- 
    -- CP-element group 1097:  join  transition  output  bypass 
    -- CP-element group 1097: predecessors 
    -- CP-element group 1097: 	1095 
    -- CP-element group 1097: 	1096 
    -- CP-element group 1097: successors 
    -- CP-element group 1097: 	1098 
    -- CP-element group 1097:  members (6) 
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/$exit
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_req
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/$exit
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/$exit
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$exit
      -- CP-element group 1097: 	 branch_block_stmt_1353/bb_36_bb_37_PhiReq/phi_stmt_2245/$exit
      -- 
    phi_stmt_2245_req_13005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2245_req_13005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1097), ack => phi_stmt_2245_req_0); -- 
    minSumDecode_cp_element_group_1097: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1097"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1095) & minSumDecode_CP_6680_elements(1096);
      gj_minSumDecode_cp_element_group_1097 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1097), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1098:  merge  place  bypass 
    -- CP-element group 1098: predecessors 
    -- CP-element group 1098: 	1089 
    -- CP-element group 1098: 	1093 
    -- CP-element group 1098: 	1097 
    -- CP-element group 1098: successors 
    -- CP-element group 1098: 	1099 
    -- CP-element group 1098:  members (1) 
      -- CP-element group 1098: 	 branch_block_stmt_1353/merge_stmt_2244_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1098) <= OrReduce(minSumDecode_CP_6680_elements(1089) & minSumDecode_CP_6680_elements(1093) & minSumDecode_CP_6680_elements(1097));
    -- CP-element group 1099:  transition  bypass 
    -- CP-element group 1099: predecessors 
    -- CP-element group 1099: 	1098 
    -- CP-element group 1099: successors 
    -- CP-element group 1099: 	1100 
    -- CP-element group 1099:  members (1) 
      -- CP-element group 1099: 	 branch_block_stmt_1353/merge_stmt_2244_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1099) <= minSumDecode_CP_6680_elements(1098);
    -- CP-element group 1100:  transition  input  no-bypass 
    -- CP-element group 1100: predecessors 
    -- CP-element group 1100: 	1099 
    -- CP-element group 1100: successors 
    -- CP-element group 1100: 	71 
    -- CP-element group 1100:  members (2) 
      -- CP-element group 1100: 	 branch_block_stmt_1353/merge_stmt_2244_PhiAck/phi_stmt_2245_ack
      -- CP-element group 1100: 	 branch_block_stmt_1353/merge_stmt_2244_PhiAck/$exit
      -- 
    phi_stmt_2245_ack_13010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2245_ack_0, ack => minSumDecode_CP_6680_elements(1100)); -- 
    -- CP-element group 1101:  fork  transition  output  bypass 
    -- CP-element group 1101: predecessors 
    -- CP-element group 1101: 	638 
    -- CP-element group 1101: successors 
    -- CP-element group 1101: 	1102 
    -- CP-element group 1101: 	1103 
    -- CP-element group 1101:  members (9) 
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Update/cr
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Update/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Sample/rr
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Sample/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/$entry
      -- CP-element group 1101: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/$entry
      -- 
    rr_13033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1101), ack => type_cast_2275_inst_req_0); -- 
    cr_13038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1101), ack => type_cast_2275_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1101) <= minSumDecode_CP_6680_elements(638);
    -- CP-element group 1102:  transition  input  no-bypass 
    -- CP-element group 1102: predecessors 
    -- CP-element group 1102: 	1101 
    -- CP-element group 1102: successors 
    -- CP-element group 1102: 	1104 
    -- CP-element group 1102:  members (2) 
      -- CP-element group 1102: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Sample/ra
      -- CP-element group 1102: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Sample/$exit
      -- 
    ra_13034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2275_inst_ack_0, ack => minSumDecode_CP_6680_elements(1102)); -- 
    -- CP-element group 1103:  transition  input  no-bypass 
    -- CP-element group 1103: predecessors 
    -- CP-element group 1103: 	1101 
    -- CP-element group 1103: successors 
    -- CP-element group 1103: 	1104 
    -- CP-element group 1103:  members (2) 
      -- CP-element group 1103: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Update/ca
      -- CP-element group 1103: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/Update/$exit
      -- 
    ca_13039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2275_inst_ack_1, ack => minSumDecode_CP_6680_elements(1103)); -- 
    -- CP-element group 1104:  join  transition  output  bypass 
    -- CP-element group 1104: predecessors 
    -- CP-element group 1104: 	1102 
    -- CP-element group 1104: 	1103 
    -- CP-element group 1104: successors 
    -- CP-element group 1104: 	1105 
    -- CP-element group 1104:  members (6) 
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_req
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/SplitProtocol/$exit
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/type_cast_2275/$exit
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/phi_stmt_2272_sources/$exit
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/phi_stmt_2272/$exit
      -- CP-element group 1104: 	 branch_block_stmt_1353/bb_37_checkIsdecodedx_xexit_PhiReq/$exit
      -- 
    phi_stmt_2272_req_13040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2272_req_13040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1104), ack => phi_stmt_2272_req_0); -- 
    minSumDecode_cp_element_group_1104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1102) & minSumDecode_CP_6680_elements(1103);
      gj_minSumDecode_cp_element_group_1104 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1105:  place  bypass 
    -- CP-element group 1105: predecessors 
    -- CP-element group 1105: 	1104 
    -- CP-element group 1105: successors 
    -- CP-element group 1105: 	1106 
    -- CP-element group 1105:  members (1) 
      -- CP-element group 1105: 	 branch_block_stmt_1353/merge_stmt_2271_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1105) <= minSumDecode_CP_6680_elements(1104);
    -- CP-element group 1106:  transition  bypass 
    -- CP-element group 1106: predecessors 
    -- CP-element group 1106: 	1105 
    -- CP-element group 1106: successors 
    -- CP-element group 1106: 	1107 
    -- CP-element group 1106:  members (1) 
      -- CP-element group 1106: 	 branch_block_stmt_1353/merge_stmt_2271_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1106) <= minSumDecode_CP_6680_elements(1105);
    -- CP-element group 1107:  transition  input  no-bypass 
    -- CP-element group 1107: predecessors 
    -- CP-element group 1107: 	1106 
    -- CP-element group 1107: successors 
    -- CP-element group 1107: 	73 
    -- CP-element group 1107:  members (2) 
      -- CP-element group 1107: 	 branch_block_stmt_1353/merge_stmt_2271_PhiAck/phi_stmt_2272_ack
      -- CP-element group 1107: 	 branch_block_stmt_1353/merge_stmt_2271_PhiAck/$exit
      -- 
    phi_stmt_2272_ack_13045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2272_ack_0, ack => minSumDecode_CP_6680_elements(1107)); -- 
    -- CP-element group 1108:  transition  bypass 
    -- CP-element group 1108: predecessors 
    -- CP-element group 1108: 	651 
    -- CP-element group 1108: successors 
    -- CP-element group 1108: 	1109 
    -- CP-element group 1108:  members (2) 
      -- CP-element group 1108: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_bb_39_PhiReq/$exit
      -- CP-element group 1108: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_bb_39_PhiReq/$entry
      -- 
    minSumDecode_CP_6680_elements(1108) <= minSumDecode_CP_6680_elements(651);
    -- CP-element group 1109:  place  bypass 
    -- CP-element group 1109: predecessors 
    -- CP-element group 1109: 	1108 
    -- CP-element group 1109: successors 
    -- CP-element group 1109: 	1110 
    -- CP-element group 1109:  members (1) 
      -- CP-element group 1109: 	 branch_block_stmt_1353/merge_stmt_2289_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1109) <= minSumDecode_CP_6680_elements(1108);
    -- CP-element group 1110:  transition  bypass 
    -- CP-element group 1110: predecessors 
    -- CP-element group 1110: 	1109 
    -- CP-element group 1110: successors 
    -- CP-element group 1110: 	75 
    -- CP-element group 1110:  members (3) 
      -- CP-element group 1110: 	 branch_block_stmt_1353/merge_stmt_2289_PhiAck/dummy
      -- CP-element group 1110: 	 branch_block_stmt_1353/merge_stmt_2289_PhiAck/$exit
      -- CP-element group 1110: 	 branch_block_stmt_1353/merge_stmt_2289_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1110) <= minSumDecode_CP_6680_elements(1109);
    -- CP-element group 1111:  transition  bypass 
    -- CP-element group 1111: predecessors 
    -- CP-element group 1111: 	665 
    -- CP-element group 1111: successors 
    -- CP-element group 1111: 	1112 
    -- CP-element group 1111:  members (2) 
      -- CP-element group 1111: 	 branch_block_stmt_1353/bb_39_bbx_xnph4x_xi_PhiReq/$exit
      -- CP-element group 1111: 	 branch_block_stmt_1353/bb_39_bbx_xnph4x_xi_PhiReq/$entry
      -- 
    minSumDecode_CP_6680_elements(1111) <= minSumDecode_CP_6680_elements(665);
    -- CP-element group 1112:  place  bypass 
    -- CP-element group 1112: predecessors 
    -- CP-element group 1112: 	1111 
    -- CP-element group 1112: successors 
    -- CP-element group 1112: 	1113 
    -- CP-element group 1112:  members (1) 
      -- CP-element group 1112: 	 branch_block_stmt_1353/merge_stmt_2305_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1112) <= minSumDecode_CP_6680_elements(1111);
    -- CP-element group 1113:  transition  bypass 
    -- CP-element group 1113: predecessors 
    -- CP-element group 1113: 	1112 
    -- CP-element group 1113: successors 
    -- CP-element group 1113: 	77 
    -- CP-element group 1113:  members (3) 
      -- CP-element group 1113: 	 branch_block_stmt_1353/merge_stmt_2305_PhiAck/dummy
      -- CP-element group 1113: 	 branch_block_stmt_1353/merge_stmt_2305_PhiAck/$exit
      -- CP-element group 1113: 	 branch_block_stmt_1353/merge_stmt_2305_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1113) <= minSumDecode_CP_6680_elements(1112);
    -- CP-element group 1114:  transition  bypass 
    -- CP-element group 1114: predecessors 
    -- CP-element group 1114: 	78 
    -- CP-element group 1114: successors 
    -- CP-element group 1114: 	1115 
    -- CP-element group 1114:  members (3) 
      -- CP-element group 1114: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/$entry
      -- CP-element group 1114: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/$entry
      -- CP-element group 1114: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/$entry
      -- 
    minSumDecode_CP_6680_elements(1114) <= minSumDecode_CP_6680_elements(78);
    -- CP-element group 1115:  transition  bypass 
    -- CP-element group 1115: predecessors 
    -- CP-element group 1115: 	1114 
    -- CP-element group 1115: successors 
    -- CP-element group 1115: 	1116 
    -- CP-element group 1115:  members (1) 
      -- CP-element group 1115: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2373_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1115) is a control-delay.
    cp_element_1115_delay: control_delay_element  generic map(name => " 1115_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1114), ack => minSumDecode_CP_6680_elements(1115), clk => clk, reset =>reset);
    -- CP-element group 1116:  transition  output  bypass 
    -- CP-element group 1116: predecessors 
    -- CP-element group 1116: 	1115 
    -- CP-element group 1116: successors 
    -- CP-element group 1116: 	1121 
    -- CP-element group 1116:  members (4) 
      -- CP-element group 1116: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/$exit
      -- CP-element group 1116: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/$exit
      -- CP-element group 1116: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/$exit
      -- CP-element group 1116: 	 branch_block_stmt_1353/bbx_xnph4x_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_req
      -- 
    phi_stmt_2369_req_13080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2369_req_13080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1116), ack => phi_stmt_2369_req_0); -- 
    minSumDecode_CP_6680_elements(1116) <= minSumDecode_CP_6680_elements(1115);
    -- CP-element group 1117:  fork  transition  output  bypass 
    -- CP-element group 1117: predecessors 
    -- CP-element group 1117: 	800 
    -- CP-element group 1117: successors 
    -- CP-element group 1117: 	1118 
    -- CP-element group 1117: 	1119 
    -- CP-element group 1117:  members (9) 
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Sample/rr
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Update/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/$entry
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Update/cr
      -- CP-element group 1117: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Sample/$entry
      -- 
    rr_13099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1117), ack => type_cast_2375_inst_req_0); -- 
    cr_13104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1117), ack => type_cast_2375_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1117) <= minSumDecode_CP_6680_elements(800);
    -- CP-element group 1118:  transition  input  no-bypass 
    -- CP-element group 1118: predecessors 
    -- CP-element group 1118: 	1117 
    -- CP-element group 1118: successors 
    -- CP-element group 1118: 	1120 
    -- CP-element group 1118:  members (2) 
      -- CP-element group 1118: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Sample/ra
      -- CP-element group 1118: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Sample/$exit
      -- 
    ra_13100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_0, ack => minSumDecode_CP_6680_elements(1118)); -- 
    -- CP-element group 1119:  transition  input  no-bypass 
    -- CP-element group 1119: predecessors 
    -- CP-element group 1119: 	1117 
    -- CP-element group 1119: successors 
    -- CP-element group 1119: 	1120 
    -- CP-element group 1119:  members (2) 
      -- CP-element group 1119: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Update/ca
      -- CP-element group 1119: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/Update/$exit
      -- 
    ca_13105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_1, ack => minSumDecode_CP_6680_elements(1119)); -- 
    -- CP-element group 1120:  join  transition  output  bypass 
    -- CP-element group 1120: predecessors 
    -- CP-element group 1120: 	1118 
    -- CP-element group 1120: 	1119 
    -- CP-element group 1120: successors 
    -- CP-element group 1120: 	1121 
    -- CP-element group 1120:  members (6) 
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_req
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/$exit
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/$exit
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/$exit
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/$exit
      -- CP-element group 1120: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_bb_41_PhiReq/phi_stmt_2369/phi_stmt_2369_sources/type_cast_2375/SplitProtocol/$exit
      -- 
    phi_stmt_2369_req_13106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2369_req_13106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1120), ack => phi_stmt_2369_req_1); -- 
    minSumDecode_cp_element_group_1120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1118) & minSumDecode_CP_6680_elements(1119);
      gj_minSumDecode_cp_element_group_1120 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1121:  merge  place  bypass 
    -- CP-element group 1121: predecessors 
    -- CP-element group 1121: 	1116 
    -- CP-element group 1121: 	1120 
    -- CP-element group 1121: successors 
    -- CP-element group 1121: 	1122 
    -- CP-element group 1121:  members (1) 
      -- CP-element group 1121: 	 branch_block_stmt_1353/merge_stmt_2368_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1121) <= OrReduce(minSumDecode_CP_6680_elements(1116) & minSumDecode_CP_6680_elements(1120));
    -- CP-element group 1122:  transition  bypass 
    -- CP-element group 1122: predecessors 
    -- CP-element group 1122: 	1121 
    -- CP-element group 1122: successors 
    -- CP-element group 1122: 	1123 
    -- CP-element group 1122:  members (1) 
      -- CP-element group 1122: 	 branch_block_stmt_1353/merge_stmt_2368_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1122) <= minSumDecode_CP_6680_elements(1121);
    -- CP-element group 1123:  transition  input  no-bypass 
    -- CP-element group 1123: predecessors 
    -- CP-element group 1123: 	1122 
    -- CP-element group 1123: successors 
    -- CP-element group 1123: 	79 
    -- CP-element group 1123:  members (2) 
      -- CP-element group 1123: 	 branch_block_stmt_1353/merge_stmt_2368_PhiAck/phi_stmt_2369_ack
      -- CP-element group 1123: 	 branch_block_stmt_1353/merge_stmt_2368_PhiAck/$exit
      -- 
    phi_stmt_2369_ack_13111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2369_ack_0, ack => minSumDecode_CP_6680_elements(1123)); -- 
    -- CP-element group 1124:  transition  bypass 
    -- CP-element group 1124: predecessors 
    -- CP-element group 1124: 	712 
    -- CP-element group 1124: successors 
    -- CP-element group 1124: 	1125 
    -- CP-element group 1124:  members (2) 
      -- CP-element group 1124: 	 branch_block_stmt_1353/bb_41_bb_42_PhiReq/$exit
      -- CP-element group 1124: 	 branch_block_stmt_1353/bb_41_bb_42_PhiReq/$entry
      -- 
    minSumDecode_CP_6680_elements(1124) <= minSumDecode_CP_6680_elements(712);
    -- CP-element group 1125:  place  bypass 
    -- CP-element group 1125: predecessors 
    -- CP-element group 1125: 	1124 
    -- CP-element group 1125: successors 
    -- CP-element group 1125: 	1126 
    -- CP-element group 1125:  members (1) 
      -- CP-element group 1125: 	 branch_block_stmt_1353/merge_stmt_2412_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1125) <= minSumDecode_CP_6680_elements(1124);
    -- CP-element group 1126:  transition  bypass 
    -- CP-element group 1126: predecessors 
    -- CP-element group 1126: 	1125 
    -- CP-element group 1126: successors 
    -- CP-element group 1126: 	81 
    -- CP-element group 1126:  members (3) 
      -- CP-element group 1126: 	 branch_block_stmt_1353/merge_stmt_2412_PhiAck/dummy
      -- CP-element group 1126: 	 branch_block_stmt_1353/merge_stmt_2412_PhiAck/$entry
      -- CP-element group 1126: 	 branch_block_stmt_1353/merge_stmt_2412_PhiAck/$exit
      -- 
    minSumDecode_CP_6680_elements(1126) <= minSumDecode_CP_6680_elements(1125);
    -- CP-element group 1127:  transition  bypass 
    -- CP-element group 1127: predecessors 
    -- CP-element group 1127: 	713 
    -- CP-element group 1127: successors 
    -- CP-element group 1127: 	1128 
    -- CP-element group 1127:  members (2) 
      -- CP-element group 1127: 	 branch_block_stmt_1353/bb_41_bb_43_PhiReq/$entry
      -- CP-element group 1127: 	 branch_block_stmt_1353/bb_41_bb_43_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1127) <= minSumDecode_CP_6680_elements(713);
    -- CP-element group 1128:  place  bypass 
    -- CP-element group 1128: predecessors 
    -- CP-element group 1128: 	1127 
    -- CP-element group 1128: successors 
    -- CP-element group 1128: 	1129 
    -- CP-element group 1128:  members (1) 
      -- CP-element group 1128: 	 branch_block_stmt_1353/merge_stmt_2423_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1128) <= minSumDecode_CP_6680_elements(1127);
    -- CP-element group 1129:  transition  bypass 
    -- CP-element group 1129: predecessors 
    -- CP-element group 1129: 	1128 
    -- CP-element group 1129: successors 
    -- CP-element group 1129: 	83 
    -- CP-element group 1129:  members (3) 
      -- CP-element group 1129: 	 branch_block_stmt_1353/merge_stmt_2423_PhiAck/dummy
      -- CP-element group 1129: 	 branch_block_stmt_1353/merge_stmt_2423_PhiAck/$entry
      -- CP-element group 1129: 	 branch_block_stmt_1353/merge_stmt_2423_PhiAck/$exit
      -- 
    minSumDecode_CP_6680_elements(1129) <= minSumDecode_CP_6680_elements(1128);
    -- CP-element group 1130:  fork  transition  output  bypass 
    -- CP-element group 1130: predecessors 
    -- CP-element group 1130: 	82 
    -- CP-element group 1130: successors 
    -- CP-element group 1130: 	1131 
    -- CP-element group 1130: 	1132 
    -- CP-element group 1130: 	1134 
    -- CP-element group 1130: 	1135 
    -- CP-element group 1130:  members (17) 
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Sample/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Sample/rr
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Update/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Update/cr
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/rr
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/$entry
      -- CP-element group 1130: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/cr
      -- 
    rr_13150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1130), ack => type_cast_2442_inst_req_0); -- 
    cr_13155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1130), ack => type_cast_2442_inst_req_1); -- 
    rr_13173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1130), ack => type_cast_2448_inst_req_0); -- 
    cr_13178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1130), ack => type_cast_2448_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1130) <= minSumDecode_CP_6680_elements(82);
    -- CP-element group 1131:  transition  input  no-bypass 
    -- CP-element group 1131: predecessors 
    -- CP-element group 1131: 	1130 
    -- CP-element group 1131: successors 
    -- CP-element group 1131: 	1133 
    -- CP-element group 1131:  members (2) 
      -- CP-element group 1131: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Sample/$exit
      -- CP-element group 1131: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Sample/ra
      -- 
    ra_13151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_0, ack => minSumDecode_CP_6680_elements(1131)); -- 
    -- CP-element group 1132:  transition  input  no-bypass 
    -- CP-element group 1132: predecessors 
    -- CP-element group 1132: 	1130 
    -- CP-element group 1132: successors 
    -- CP-element group 1132: 	1133 
    -- CP-element group 1132:  members (2) 
      -- CP-element group 1132: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Update/$exit
      -- CP-element group 1132: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/Update/ca
      -- 
    ca_13156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_1, ack => minSumDecode_CP_6680_elements(1132)); -- 
    -- CP-element group 1133:  join  transition  output  bypass 
    -- CP-element group 1133: predecessors 
    -- CP-element group 1133: 	1131 
    -- CP-element group 1133: 	1132 
    -- CP-element group 1133: successors 
    -- CP-element group 1133: 	1137 
    -- CP-element group 1133:  members (5) 
      -- CP-element group 1133: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/SplitProtocol/$exit
      -- CP-element group 1133: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2442/$exit
      -- CP-element group 1133: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/$exit
      -- CP-element group 1133: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/$exit
      -- CP-element group 1133: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_req
      -- 
    phi_stmt_2439_req_13157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2439_req_13157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1133), ack => phi_stmt_2439_req_0); -- 
    minSumDecode_cp_element_group_1133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1131) & minSumDecode_CP_6680_elements(1132);
      gj_minSumDecode_cp_element_group_1133 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1134:  transition  input  no-bypass 
    -- CP-element group 1134: predecessors 
    -- CP-element group 1134: 	1130 
    -- CP-element group 1134: successors 
    -- CP-element group 1134: 	1136 
    -- CP-element group 1134:  members (2) 
      -- CP-element group 1134: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/$exit
      -- CP-element group 1134: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/ra
      -- 
    ra_13174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_0, ack => minSumDecode_CP_6680_elements(1134)); -- 
    -- CP-element group 1135:  transition  input  no-bypass 
    -- CP-element group 1135: predecessors 
    -- CP-element group 1135: 	1130 
    -- CP-element group 1135: successors 
    -- CP-element group 1135: 	1136 
    -- CP-element group 1135:  members (2) 
      -- CP-element group 1135: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/$exit
      -- CP-element group 1135: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/ca
      -- 
    ca_13179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_1, ack => minSumDecode_CP_6680_elements(1135)); -- 
    -- CP-element group 1136:  join  transition  output  bypass 
    -- CP-element group 1136: predecessors 
    -- CP-element group 1136: 	1134 
    -- CP-element group 1136: 	1135 
    -- CP-element group 1136: successors 
    -- CP-element group 1136: 	1137 
    -- CP-element group 1136:  members (5) 
      -- CP-element group 1136: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/$exit
      -- CP-element group 1136: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$exit
      -- CP-element group 1136: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/$exit
      -- CP-element group 1136: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/$exit
      -- CP-element group 1136: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_req
      -- 
    phi_stmt_2445_req_13180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2445_req_13180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1136), ack => phi_stmt_2445_req_0); -- 
    minSumDecode_cp_element_group_1136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1134) & minSumDecode_CP_6680_elements(1135);
      gj_minSumDecode_cp_element_group_1136 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1137:  join  transition  bypass 
    -- CP-element group 1137: predecessors 
    -- CP-element group 1137: 	1133 
    -- CP-element group 1137: 	1136 
    -- CP-element group 1137: successors 
    -- CP-element group 1137: 	1146 
    -- CP-element group 1137:  members (1) 
      -- CP-element group 1137: 	 branch_block_stmt_1353/bb_42_bb_44_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1133) & minSumDecode_CP_6680_elements(1136);
      gj_minSumDecode_cp_element_group_1137 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1138:  fork  transition  output  bypass 
    -- CP-element group 1138: predecessors 
    -- CP-element group 1138: 	84 
    -- CP-element group 1138: successors 
    -- CP-element group 1138: 	1139 
    -- CP-element group 1138: 	1140 
    -- CP-element group 1138: 	1142 
    -- CP-element group 1138: 	1143 
    -- CP-element group 1138:  members (17) 
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Sample/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Sample/rr
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Update/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Update/cr
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/rr
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/$entry
      -- CP-element group 1138: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/cr
      -- 
    rr_13199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1138), ack => type_cast_2444_inst_req_0); -- 
    cr_13204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1138), ack => type_cast_2444_inst_req_1); -- 
    rr_13222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1138), ack => type_cast_2450_inst_req_0); -- 
    cr_13227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1138), ack => type_cast_2450_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1138) <= minSumDecode_CP_6680_elements(84);
    -- CP-element group 1139:  transition  input  no-bypass 
    -- CP-element group 1139: predecessors 
    -- CP-element group 1139: 	1138 
    -- CP-element group 1139: successors 
    -- CP-element group 1139: 	1141 
    -- CP-element group 1139:  members (2) 
      -- CP-element group 1139: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Sample/$exit
      -- CP-element group 1139: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Sample/ra
      -- 
    ra_13200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_0, ack => minSumDecode_CP_6680_elements(1139)); -- 
    -- CP-element group 1140:  transition  input  no-bypass 
    -- CP-element group 1140: predecessors 
    -- CP-element group 1140: 	1138 
    -- CP-element group 1140: successors 
    -- CP-element group 1140: 	1141 
    -- CP-element group 1140:  members (2) 
      -- CP-element group 1140: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Update/$exit
      -- CP-element group 1140: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/Update/ca
      -- 
    ca_13205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_1, ack => minSumDecode_CP_6680_elements(1140)); -- 
    -- CP-element group 1141:  join  transition  output  bypass 
    -- CP-element group 1141: predecessors 
    -- CP-element group 1141: 	1139 
    -- CP-element group 1141: 	1140 
    -- CP-element group 1141: successors 
    -- CP-element group 1141: 	1145 
    -- CP-element group 1141:  members (5) 
      -- CP-element group 1141: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/$exit
      -- CP-element group 1141: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/$exit
      -- CP-element group 1141: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/$exit
      -- CP-element group 1141: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_sources/type_cast_2444/SplitProtocol/$exit
      -- CP-element group 1141: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2439/phi_stmt_2439_req
      -- 
    phi_stmt_2439_req_13206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2439_req_13206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1141), ack => phi_stmt_2439_req_1); -- 
    minSumDecode_cp_element_group_1141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1139) & minSumDecode_CP_6680_elements(1140);
      gj_minSumDecode_cp_element_group_1141 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1142:  transition  input  no-bypass 
    -- CP-element group 1142: predecessors 
    -- CP-element group 1142: 	1138 
    -- CP-element group 1142: successors 
    -- CP-element group 1142: 	1144 
    -- CP-element group 1142:  members (2) 
      -- CP-element group 1142: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/$exit
      -- CP-element group 1142: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/ra
      -- 
    ra_13223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_0, ack => minSumDecode_CP_6680_elements(1142)); -- 
    -- CP-element group 1143:  transition  input  no-bypass 
    -- CP-element group 1143: predecessors 
    -- CP-element group 1143: 	1138 
    -- CP-element group 1143: successors 
    -- CP-element group 1143: 	1144 
    -- CP-element group 1143:  members (2) 
      -- CP-element group 1143: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/$exit
      -- CP-element group 1143: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/ca
      -- 
    ca_13228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_1, ack => minSumDecode_CP_6680_elements(1143)); -- 
    -- CP-element group 1144:  join  transition  output  bypass 
    -- CP-element group 1144: predecessors 
    -- CP-element group 1144: 	1142 
    -- CP-element group 1144: 	1143 
    -- CP-element group 1144: successors 
    -- CP-element group 1144: 	1145 
    -- CP-element group 1144:  members (5) 
      -- CP-element group 1144: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/$exit
      -- CP-element group 1144: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$exit
      -- CP-element group 1144: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/$exit
      -- CP-element group 1144: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/$exit
      -- CP-element group 1144: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/phi_stmt_2445/phi_stmt_2445_req
      -- 
    phi_stmt_2445_req_13229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2445_req_13229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1144), ack => phi_stmt_2445_req_1); -- 
    minSumDecode_cp_element_group_1144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1142) & minSumDecode_CP_6680_elements(1143);
      gj_minSumDecode_cp_element_group_1144 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1145:  join  transition  bypass 
    -- CP-element group 1145: predecessors 
    -- CP-element group 1145: 	1141 
    -- CP-element group 1145: 	1144 
    -- CP-element group 1145: successors 
    -- CP-element group 1145: 	1146 
    -- CP-element group 1145:  members (1) 
      -- CP-element group 1145: 	 branch_block_stmt_1353/bb_43_bb_44_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1141) & minSumDecode_CP_6680_elements(1144);
      gj_minSumDecode_cp_element_group_1145 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1146:  merge  place  bypass 
    -- CP-element group 1146: predecessors 
    -- CP-element group 1146: 	1137 
    -- CP-element group 1146: 	1145 
    -- CP-element group 1146: successors 
    -- CP-element group 1146: 	1147 
    -- CP-element group 1146:  members (1) 
      -- CP-element group 1146: 	 branch_block_stmt_1353/merge_stmt_2438_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1146) <= OrReduce(minSumDecode_CP_6680_elements(1137) & minSumDecode_CP_6680_elements(1145));
    -- CP-element group 1147:  fork  transition  bypass 
    -- CP-element group 1147: predecessors 
    -- CP-element group 1147: 	1146 
    -- CP-element group 1147: successors 
    -- CP-element group 1147: 	1148 
    -- CP-element group 1147: 	1149 
    -- CP-element group 1147:  members (1) 
      -- CP-element group 1147: 	 branch_block_stmt_1353/merge_stmt_2438_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1147) <= minSumDecode_CP_6680_elements(1146);
    -- CP-element group 1148:  transition  input  no-bypass 
    -- CP-element group 1148: predecessors 
    -- CP-element group 1148: 	1147 
    -- CP-element group 1148: successors 
    -- CP-element group 1148: 	1150 
    -- CP-element group 1148:  members (1) 
      -- CP-element group 1148: 	 branch_block_stmt_1353/merge_stmt_2438_PhiAck/phi_stmt_2439_ack
      -- 
    phi_stmt_2439_ack_13234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2439_ack_0, ack => minSumDecode_CP_6680_elements(1148)); -- 
    -- CP-element group 1149:  transition  input  no-bypass 
    -- CP-element group 1149: predecessors 
    -- CP-element group 1149: 	1147 
    -- CP-element group 1149: successors 
    -- CP-element group 1149: 	1150 
    -- CP-element group 1149:  members (1) 
      -- CP-element group 1149: 	 branch_block_stmt_1353/merge_stmt_2438_PhiAck/phi_stmt_2445_ack
      -- 
    phi_stmt_2445_ack_13235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2445_ack_0, ack => minSumDecode_CP_6680_elements(1149)); -- 
    -- CP-element group 1150:  join  transition  bypass 
    -- CP-element group 1150: predecessors 
    -- CP-element group 1150: 	1148 
    -- CP-element group 1150: 	1149 
    -- CP-element group 1150: successors 
    -- CP-element group 1150: 	85 
    -- CP-element group 1150:  members (1) 
      -- CP-element group 1150: 	 branch_block_stmt_1353/merge_stmt_2438_PhiAck/$exit
      -- 
    minSumDecode_cp_element_group_1150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1148) & minSumDecode_CP_6680_elements(1149);
      gj_minSumDecode_cp_element_group_1150 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1151:  transition  bypass 
    -- CP-element group 1151: predecessors 
    -- CP-element group 1151: 	738 
    -- CP-element group 1151: successors 
    -- CP-element group 1151: 	1152 
    -- CP-element group 1151:  members (2) 
      -- CP-element group 1151: 	 branch_block_stmt_1353/bb_44_bbx_xnphx_xi36_PhiReq/$entry
      -- CP-element group 1151: 	 branch_block_stmt_1353/bb_44_bbx_xnphx_xi36_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1151) <= minSumDecode_CP_6680_elements(738);
    -- CP-element group 1152:  place  bypass 
    -- CP-element group 1152: predecessors 
    -- CP-element group 1152: 	1151 
    -- CP-element group 1152: successors 
    -- CP-element group 1152: 	1153 
    -- CP-element group 1152:  members (1) 
      -- CP-element group 1152: 	 branch_block_stmt_1353/merge_stmt_2464_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1152) <= minSumDecode_CP_6680_elements(1151);
    -- CP-element group 1153:  transition  bypass 
    -- CP-element group 1153: predecessors 
    -- CP-element group 1153: 	1152 
    -- CP-element group 1153: successors 
    -- CP-element group 1153: 	87 
    -- CP-element group 1153:  members (3) 
      -- CP-element group 1153: 	 branch_block_stmt_1353/merge_stmt_2464_PhiAck/$entry
      -- CP-element group 1153: 	 branch_block_stmt_1353/merge_stmt_2464_PhiAck/$exit
      -- CP-element group 1153: 	 branch_block_stmt_1353/merge_stmt_2464_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1153) <= minSumDecode_CP_6680_elements(1152);
    -- CP-element group 1154:  fork  transition  output  bypass 
    -- CP-element group 1154: predecessors 
    -- CP-element group 1154: 	786 
    -- CP-element group 1154: successors 
    -- CP-element group 1154: 	1155 
    -- CP-element group 1154: 	1156 
    -- CP-element group 1154:  members (9) 
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Sample/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Sample/rr
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Update/$entry
      -- CP-element group 1154: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Update/cr
      -- 
    rr_13266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1154), ack => type_cast_2479_inst_req_0); -- 
    cr_13271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1154), ack => type_cast_2479_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1154) <= minSumDecode_CP_6680_elements(786);
    -- CP-element group 1155:  transition  input  no-bypass 
    -- CP-element group 1155: predecessors 
    -- CP-element group 1155: 	1154 
    -- CP-element group 1155: successors 
    -- CP-element group 1155: 	1157 
    -- CP-element group 1155:  members (2) 
      -- CP-element group 1155: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Sample/$exit
      -- CP-element group 1155: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Sample/ra
      -- 
    ra_13267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2479_inst_ack_0, ack => minSumDecode_CP_6680_elements(1155)); -- 
    -- CP-element group 1156:  transition  input  no-bypass 
    -- CP-element group 1156: predecessors 
    -- CP-element group 1156: 	1154 
    -- CP-element group 1156: successors 
    -- CP-element group 1156: 	1157 
    -- CP-element group 1156:  members (2) 
      -- CP-element group 1156: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Update/$exit
      -- CP-element group 1156: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/Update/ca
      -- 
    ca_13272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2479_inst_ack_1, ack => minSumDecode_CP_6680_elements(1156)); -- 
    -- CP-element group 1157:  join  transition  output  bypass 
    -- CP-element group 1157: predecessors 
    -- CP-element group 1157: 	1155 
    -- CP-element group 1157: 	1156 
    -- CP-element group 1157: successors 
    -- CP-element group 1157: 	1161 
    -- CP-element group 1157:  members (6) 
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/$exit
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/$exit
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/$exit
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/$exit
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2479/SplitProtocol/$exit
      -- CP-element group 1157: 	 branch_block_stmt_1353/bb_46_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_req
      -- 
    phi_stmt_2473_req_13273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2473_req_13273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1157), ack => phi_stmt_2473_req_1); -- 
    minSumDecode_cp_element_group_1157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1155) & minSumDecode_CP_6680_elements(1156);
      gj_minSumDecode_cp_element_group_1157 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1158:  transition  bypass 
    -- CP-element group 1158: predecessors 
    -- CP-element group 1158: 	88 
    -- CP-element group 1158: successors 
    -- CP-element group 1158: 	1159 
    -- CP-element group 1158:  members (3) 
      -- CP-element group 1158: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/$entry
      -- CP-element group 1158: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/$entry
      -- CP-element group 1158: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1158) <= minSumDecode_CP_6680_elements(88);
    -- CP-element group 1159:  transition  bypass 
    -- CP-element group 1159: predecessors 
    -- CP-element group 1159: 	1158 
    -- CP-element group 1159: successors 
    -- CP-element group 1159: 	1160 
    -- CP-element group 1159:  members (1) 
      -- CP-element group 1159: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/type_cast_2477_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1159) is a control-delay.
    cp_element_1159_delay: control_delay_element  generic map(name => " 1159_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1158), ack => minSumDecode_CP_6680_elements(1159), clk => clk, reset =>reset);
    -- CP-element group 1160:  transition  output  bypass 
    -- CP-element group 1160: predecessors 
    -- CP-element group 1160: 	1159 
    -- CP-element group 1160: successors 
    -- CP-element group 1160: 	1161 
    -- CP-element group 1160:  members (4) 
      -- CP-element group 1160: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/$exit
      -- CP-element group 1160: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/$exit
      -- CP-element group 1160: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_sources/$exit
      -- CP-element group 1160: 	 branch_block_stmt_1353/bbx_xnphx_xi36_bb_46_PhiReq/phi_stmt_2473/phi_stmt_2473_req
      -- 
    phi_stmt_2473_req_13284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2473_req_13284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1160), ack => phi_stmt_2473_req_0); -- 
    minSumDecode_CP_6680_elements(1160) <= minSumDecode_CP_6680_elements(1159);
    -- CP-element group 1161:  merge  place  bypass 
    -- CP-element group 1161: predecessors 
    -- CP-element group 1161: 	1157 
    -- CP-element group 1161: 	1160 
    -- CP-element group 1161: successors 
    -- CP-element group 1161: 	1162 
    -- CP-element group 1161:  members (1) 
      -- CP-element group 1161: 	 branch_block_stmt_1353/merge_stmt_2472_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1161) <= OrReduce(minSumDecode_CP_6680_elements(1157) & minSumDecode_CP_6680_elements(1160));
    -- CP-element group 1162:  transition  bypass 
    -- CP-element group 1162: predecessors 
    -- CP-element group 1162: 	1161 
    -- CP-element group 1162: successors 
    -- CP-element group 1162: 	1163 
    -- CP-element group 1162:  members (1) 
      -- CP-element group 1162: 	 branch_block_stmt_1353/merge_stmt_2472_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1162) <= minSumDecode_CP_6680_elements(1161);
    -- CP-element group 1163:  transition  input  no-bypass 
    -- CP-element group 1163: predecessors 
    -- CP-element group 1163: 	1162 
    -- CP-element group 1163: successors 
    -- CP-element group 1163: 	89 
    -- CP-element group 1163:  members (2) 
      -- CP-element group 1163: 	 branch_block_stmt_1353/merge_stmt_2472_PhiAck/$exit
      -- CP-element group 1163: 	 branch_block_stmt_1353/merge_stmt_2472_PhiAck/phi_stmt_2473_ack
      -- 
    phi_stmt_2473_ack_13289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2473_ack_0, ack => minSumDecode_CP_6680_elements(1163)); -- 
    -- CP-element group 1164:  transition  bypass 
    -- CP-element group 1164: predecessors 
    -- CP-element group 1164: 	785 
    -- CP-element group 1164: successors 
    -- CP-element group 1164: 	1165 
    -- CP-element group 1164:  members (2) 
      -- CP-element group 1164: 	 branch_block_stmt_1353/bb_46_xx_x_crit_edgex_xix_xloopexit_PhiReq/$entry
      -- CP-element group 1164: 	 branch_block_stmt_1353/bb_46_xx_x_crit_edgex_xix_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1164) <= minSumDecode_CP_6680_elements(785);
    -- CP-element group 1165:  place  bypass 
    -- CP-element group 1165: predecessors 
    -- CP-element group 1165: 	1164 
    -- CP-element group 1165: successors 
    -- CP-element group 1165: 	1166 
    -- CP-element group 1165:  members (1) 
      -- CP-element group 1165: 	 branch_block_stmt_1353/merge_stmt_2564_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1165) <= minSumDecode_CP_6680_elements(1164);
    -- CP-element group 1166:  transition  bypass 
    -- CP-element group 1166: predecessors 
    -- CP-element group 1166: 	1165 
    -- CP-element group 1166: successors 
    -- CP-element group 1166: 	91 
    -- CP-element group 1166:  members (3) 
      -- CP-element group 1166: 	 branch_block_stmt_1353/merge_stmt_2564_PhiAck/$entry
      -- CP-element group 1166: 	 branch_block_stmt_1353/merge_stmt_2564_PhiAck/$exit
      -- CP-element group 1166: 	 branch_block_stmt_1353/merge_stmt_2564_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1166) <= minSumDecode_CP_6680_elements(1165);
    -- CP-element group 1167:  transition  bypass 
    -- CP-element group 1167: predecessors 
    -- CP-element group 1167: 	737 
    -- CP-element group 1167: successors 
    -- CP-element group 1167: 	1169 
    -- CP-element group 1167:  members (2) 
      -- CP-element group 1167: 	 branch_block_stmt_1353/bb_44_xx_x_crit_edgex_xi_PhiReq/$entry
      -- CP-element group 1167: 	 branch_block_stmt_1353/bb_44_xx_x_crit_edgex_xi_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1167) <= minSumDecode_CP_6680_elements(737);
    -- CP-element group 1168:  transition  bypass 
    -- CP-element group 1168: predecessors 
    -- CP-element group 1168: 	91 
    -- CP-element group 1168: successors 
    -- CP-element group 1168: 	1169 
    -- CP-element group 1168:  members (2) 
      -- CP-element group 1168: 	 branch_block_stmt_1353/xx_x_crit_edgex_xix_xloopexit_xx_x_crit_edgex_xi_PhiReq/$entry
      -- CP-element group 1168: 	 branch_block_stmt_1353/xx_x_crit_edgex_xix_xloopexit_xx_x_crit_edgex_xi_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1168) <= minSumDecode_CP_6680_elements(91);
    -- CP-element group 1169:  merge  place  bypass 
    -- CP-element group 1169: predecessors 
    -- CP-element group 1169: 	1167 
    -- CP-element group 1169: 	1168 
    -- CP-element group 1169: successors 
    -- CP-element group 1169: 	1170 
    -- CP-element group 1169:  members (1) 
      -- CP-element group 1169: 	 branch_block_stmt_1353/merge_stmt_2566_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1169) <= OrReduce(minSumDecode_CP_6680_elements(1167) & minSumDecode_CP_6680_elements(1168));
    -- CP-element group 1170:  transition  bypass 
    -- CP-element group 1170: predecessors 
    -- CP-element group 1170: 	1169 
    -- CP-element group 1170: successors 
    -- CP-element group 1170: 	92 
    -- CP-element group 1170:  members (3) 
      -- CP-element group 1170: 	 branch_block_stmt_1353/merge_stmt_2566_PhiAck/$entry
      -- CP-element group 1170: 	 branch_block_stmt_1353/merge_stmt_2566_PhiAck/$exit
      -- CP-element group 1170: 	 branch_block_stmt_1353/merge_stmt_2566_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1170) <= minSumDecode_CP_6680_elements(1169);
    -- CP-element group 1171:  transition  bypass 
    -- CP-element group 1171: predecessors 
    -- CP-element group 1171: 	799 
    -- CP-element group 1171: successors 
    -- CP-element group 1171: 	1172 
    -- CP-element group 1171:  members (2) 
      -- CP-element group 1171: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_updateMessagex_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 1171: 	 branch_block_stmt_1353/xx_x_crit_edgex_xi_updateMessagex_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1171) <= minSumDecode_CP_6680_elements(799);
    -- CP-element group 1172:  place  bypass 
    -- CP-element group 1172: predecessors 
    -- CP-element group 1172: 	1171 
    -- CP-element group 1172: successors 
    -- CP-element group 1172: 	1173 
    -- CP-element group 1172:  members (1) 
      -- CP-element group 1172: 	 branch_block_stmt_1353/merge_stmt_2584_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1172) <= minSumDecode_CP_6680_elements(1171);
    -- CP-element group 1173:  transition  bypass 
    -- CP-element group 1173: predecessors 
    -- CP-element group 1173: 	1172 
    -- CP-element group 1173: successors 
    -- CP-element group 1173: 	94 
    -- CP-element group 1173:  members (3) 
      -- CP-element group 1173: 	 branch_block_stmt_1353/merge_stmt_2584_PhiAck/$entry
      -- CP-element group 1173: 	 branch_block_stmt_1353/merge_stmt_2584_PhiAck/$exit
      -- CP-element group 1173: 	 branch_block_stmt_1353/merge_stmt_2584_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1173) <= minSumDecode_CP_6680_elements(1172);
    -- CP-element group 1174:  transition  bypass 
    -- CP-element group 1174: predecessors 
    -- CP-element group 1174: 	664 
    -- CP-element group 1174: successors 
    -- CP-element group 1174: 	1176 
    -- CP-element group 1174:  members (2) 
      -- CP-element group 1174: 	 branch_block_stmt_1353/bb_39_updateMessagex_xexit_PhiReq/$entry
      -- CP-element group 1174: 	 branch_block_stmt_1353/bb_39_updateMessagex_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1174) <= minSumDecode_CP_6680_elements(664);
    -- CP-element group 1175:  transition  bypass 
    -- CP-element group 1175: predecessors 
    -- CP-element group 1175: 	94 
    -- CP-element group 1175: successors 
    -- CP-element group 1175: 	1176 
    -- CP-element group 1175:  members (2) 
      -- CP-element group 1175: 	 branch_block_stmt_1353/updateMessagex_xexitx_xloopexit_updateMessagex_xexit_PhiReq/$entry
      -- CP-element group 1175: 	 branch_block_stmt_1353/updateMessagex_xexitx_xloopexit_updateMessagex_xexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1175) <= minSumDecode_CP_6680_elements(94);
    -- CP-element group 1176:  merge  place  bypass 
    -- CP-element group 1176: predecessors 
    -- CP-element group 1176: 	1174 
    -- CP-element group 1176: 	1175 
    -- CP-element group 1176: successors 
    -- CP-element group 1176: 	1177 
    -- CP-element group 1176:  members (1) 
      -- CP-element group 1176: 	 branch_block_stmt_1353/merge_stmt_2586_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1176) <= OrReduce(minSumDecode_CP_6680_elements(1174) & minSumDecode_CP_6680_elements(1175));
    -- CP-element group 1177:  transition  bypass 
    -- CP-element group 1177: predecessors 
    -- CP-element group 1177: 	1176 
    -- CP-element group 1177: successors 
    -- CP-element group 1177: 	95 
    -- CP-element group 1177:  members (3) 
      -- CP-element group 1177: 	 branch_block_stmt_1353/merge_stmt_2586_PhiAck/$entry
      -- CP-element group 1177: 	 branch_block_stmt_1353/merge_stmt_2586_PhiAck/$exit
      -- CP-element group 1177: 	 branch_block_stmt_1353/merge_stmt_2586_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1177) <= minSumDecode_CP_6680_elements(1176);
    -- CP-element group 1178:  fork  transition  output  bypass 
    -- CP-element group 1178: predecessors 
    -- CP-element group 1178: 	650 
    -- CP-element group 1178: successors 
    -- CP-element group 1178: 	1179 
    -- CP-element group 1178: 	1180 
    -- CP-element group 1178: 	1182 
    -- CP-element group 1178: 	1183 
    -- CP-element group 1178:  members (17) 
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Sample/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Sample/rr
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Update/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Update/cr
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Sample/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Sample/rr
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Update/$entry
      -- CP-element group 1178: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Update/cr
      -- 
    rr_13354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1178), ack => type_cast_2598_inst_req_0); -- 
    cr_13359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1178), ack => type_cast_2598_inst_req_1); -- 
    rr_13377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1178), ack => type_cast_2604_inst_req_0); -- 
    cr_13382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1178), ack => type_cast_2604_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1178) <= minSumDecode_CP_6680_elements(650);
    -- CP-element group 1179:  transition  input  no-bypass 
    -- CP-element group 1179: predecessors 
    -- CP-element group 1179: 	1178 
    -- CP-element group 1179: successors 
    -- CP-element group 1179: 	1181 
    -- CP-element group 1179:  members (2) 
      -- CP-element group 1179: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Sample/$exit
      -- CP-element group 1179: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Sample/ra
      -- 
    ra_13355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_0, ack => minSumDecode_CP_6680_elements(1179)); -- 
    -- CP-element group 1180:  transition  input  no-bypass 
    -- CP-element group 1180: predecessors 
    -- CP-element group 1180: 	1178 
    -- CP-element group 1180: successors 
    -- CP-element group 1180: 	1181 
    -- CP-element group 1180:  members (2) 
      -- CP-element group 1180: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Update/$exit
      -- CP-element group 1180: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/Update/ca
      -- 
    ca_13360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_1, ack => minSumDecode_CP_6680_elements(1180)); -- 
    -- CP-element group 1181:  join  transition  output  bypass 
    -- CP-element group 1181: predecessors 
    -- CP-element group 1181: 	1179 
    -- CP-element group 1181: 	1180 
    -- CP-element group 1181: successors 
    -- CP-element group 1181: 	1185 
    -- CP-element group 1181:  members (5) 
      -- CP-element group 1181: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/$exit
      -- CP-element group 1181: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$exit
      -- CP-element group 1181: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/$exit
      -- CP-element group 1181: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2598/SplitProtocol/$exit
      -- CP-element group 1181: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_req
      -- 
    phi_stmt_2595_req_13361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2595_req_13361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1181), ack => phi_stmt_2595_req_0); -- 
    minSumDecode_cp_element_group_1181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1179) & minSumDecode_CP_6680_elements(1180);
      gj_minSumDecode_cp_element_group_1181 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1182:  transition  input  no-bypass 
    -- CP-element group 1182: predecessors 
    -- CP-element group 1182: 	1178 
    -- CP-element group 1182: successors 
    -- CP-element group 1182: 	1184 
    -- CP-element group 1182:  members (2) 
      -- CP-element group 1182: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Sample/$exit
      -- CP-element group 1182: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Sample/ra
      -- 
    ra_13378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2604_inst_ack_0, ack => minSumDecode_CP_6680_elements(1182)); -- 
    -- CP-element group 1183:  transition  input  no-bypass 
    -- CP-element group 1183: predecessors 
    -- CP-element group 1183: 	1178 
    -- CP-element group 1183: successors 
    -- CP-element group 1183: 	1184 
    -- CP-element group 1183:  members (2) 
      -- CP-element group 1183: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Update/$exit
      -- CP-element group 1183: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/Update/ca
      -- 
    ca_13383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2604_inst_ack_1, ack => minSumDecode_CP_6680_elements(1183)); -- 
    -- CP-element group 1184:  join  transition  output  bypass 
    -- CP-element group 1184: predecessors 
    -- CP-element group 1184: 	1182 
    -- CP-element group 1184: 	1183 
    -- CP-element group 1184: successors 
    -- CP-element group 1184: 	1185 
    -- CP-element group 1184:  members (5) 
      -- CP-element group 1184: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/$exit
      -- CP-element group 1184: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/$exit
      -- CP-element group 1184: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/$exit
      -- CP-element group 1184: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2604/SplitProtocol/$exit
      -- CP-element group 1184: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_req
      -- 
    phi_stmt_2601_req_13384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_req_13384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1184), ack => phi_stmt_2601_req_0); -- 
    minSumDecode_cp_element_group_1184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1182) & minSumDecode_CP_6680_elements(1183);
      gj_minSumDecode_cp_element_group_1184 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1185:  join  transition  bypass 
    -- CP-element group 1185: predecessors 
    -- CP-element group 1185: 	1181 
    -- CP-element group 1185: 	1184 
    -- CP-element group 1185: successors 
    -- CP-element group 1185: 	1194 
    -- CP-element group 1185:  members (1) 
      -- CP-element group 1185: 	 branch_block_stmt_1353/checkIsdecodedx_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1181) & minSumDecode_CP_6680_elements(1184);
      gj_minSumDecode_cp_element_group_1185 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1186:  fork  transition  output  bypass 
    -- CP-element group 1186: predecessors 
    -- CP-element group 1186: 	352 
    -- CP-element group 1186: successors 
    -- CP-element group 1186: 	1187 
    -- CP-element group 1186: 	1188 
    -- CP-element group 1186: 	1190 
    -- CP-element group 1186: 	1191 
    -- CP-element group 1186:  members (17) 
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Sample/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Sample/rr
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Update/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Update/cr
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Sample/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Sample/rr
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Update/$entry
      -- CP-element group 1186: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Update/cr
      -- 
    rr_13403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1186), ack => type_cast_2600_inst_req_0); -- 
    cr_13408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1186), ack => type_cast_2600_inst_req_1); -- 
    rr_13426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1186), ack => type_cast_2606_inst_req_0); -- 
    cr_13431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1186), ack => type_cast_2606_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1186) <= minSumDecode_CP_6680_elements(352);
    -- CP-element group 1187:  transition  input  no-bypass 
    -- CP-element group 1187: predecessors 
    -- CP-element group 1187: 	1186 
    -- CP-element group 1187: successors 
    -- CP-element group 1187: 	1189 
    -- CP-element group 1187:  members (2) 
      -- CP-element group 1187: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Sample/$exit
      -- CP-element group 1187: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Sample/ra
      -- 
    ra_13404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_0, ack => minSumDecode_CP_6680_elements(1187)); -- 
    -- CP-element group 1188:  transition  input  no-bypass 
    -- CP-element group 1188: predecessors 
    -- CP-element group 1188: 	1186 
    -- CP-element group 1188: successors 
    -- CP-element group 1188: 	1189 
    -- CP-element group 1188:  members (2) 
      -- CP-element group 1188: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Update/$exit
      -- CP-element group 1188: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/Update/ca
      -- 
    ca_13409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_1, ack => minSumDecode_CP_6680_elements(1188)); -- 
    -- CP-element group 1189:  join  transition  output  bypass 
    -- CP-element group 1189: predecessors 
    -- CP-element group 1189: 	1187 
    -- CP-element group 1189: 	1188 
    -- CP-element group 1189: successors 
    -- CP-element group 1189: 	1193 
    -- CP-element group 1189:  members (5) 
      -- CP-element group 1189: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/$exit
      -- CP-element group 1189: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/$exit
      -- CP-element group 1189: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/$exit
      -- CP-element group 1189: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_sources/type_cast_2600/SplitProtocol/$exit
      -- CP-element group 1189: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2595/phi_stmt_2595_req
      -- 
    phi_stmt_2595_req_13410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2595_req_13410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1189), ack => phi_stmt_2595_req_1); -- 
    minSumDecode_cp_element_group_1189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1187) & minSumDecode_CP_6680_elements(1188);
      gj_minSumDecode_cp_element_group_1189 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1190:  transition  input  no-bypass 
    -- CP-element group 1190: predecessors 
    -- CP-element group 1190: 	1186 
    -- CP-element group 1190: successors 
    -- CP-element group 1190: 	1192 
    -- CP-element group 1190:  members (2) 
      -- CP-element group 1190: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Sample/$exit
      -- CP-element group 1190: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Sample/ra
      -- 
    ra_13427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_0, ack => minSumDecode_CP_6680_elements(1190)); -- 
    -- CP-element group 1191:  transition  input  no-bypass 
    -- CP-element group 1191: predecessors 
    -- CP-element group 1191: 	1186 
    -- CP-element group 1191: successors 
    -- CP-element group 1191: 	1192 
    -- CP-element group 1191:  members (2) 
      -- CP-element group 1191: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Update/$exit
      -- CP-element group 1191: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/Update/ca
      -- 
    ca_13432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_1, ack => minSumDecode_CP_6680_elements(1191)); -- 
    -- CP-element group 1192:  join  transition  output  bypass 
    -- CP-element group 1192: predecessors 
    -- CP-element group 1192: 	1190 
    -- CP-element group 1192: 	1191 
    -- CP-element group 1192: successors 
    -- CP-element group 1192: 	1193 
    -- CP-element group 1192:  members (5) 
      -- CP-element group 1192: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/$exit
      -- CP-element group 1192: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/$exit
      -- CP-element group 1192: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/$exit
      -- CP-element group 1192: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_sources/type_cast_2606/SplitProtocol/$exit
      -- CP-element group 1192: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/phi_stmt_2601/phi_stmt_2601_req
      -- 
    phi_stmt_2601_req_13433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_req_13433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1192), ack => phi_stmt_2601_req_1); -- 
    minSumDecode_cp_element_group_1192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1190) & minSumDecode_CP_6680_elements(1191);
      gj_minSumDecode_cp_element_group_1192 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1193:  join  transition  bypass 
    -- CP-element group 1193: predecessors 
    -- CP-element group 1193: 	1189 
    -- CP-element group 1193: 	1192 
    -- CP-element group 1193: successors 
    -- CP-element group 1193: 	1194 
    -- CP-element group 1193:  members (1) 
      -- CP-element group 1193: 	 branch_block_stmt_1353/initializeMessagex_xexit_checkIsdecodedx_xexitx_xthread_PhiReq/$exit
      -- 
    minSumDecode_cp_element_group_1193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1189) & minSumDecode_CP_6680_elements(1192);
      gj_minSumDecode_cp_element_group_1193 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1194:  merge  place  bypass 
    -- CP-element group 1194: predecessors 
    -- CP-element group 1194: 	1185 
    -- CP-element group 1194: 	1193 
    -- CP-element group 1194: successors 
    -- CP-element group 1194: 	1195 
    -- CP-element group 1194:  members (1) 
      -- CP-element group 1194: 	 branch_block_stmt_1353/merge_stmt_2594_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1194) <= OrReduce(minSumDecode_CP_6680_elements(1185) & minSumDecode_CP_6680_elements(1193));
    -- CP-element group 1195:  fork  transition  bypass 
    -- CP-element group 1195: predecessors 
    -- CP-element group 1195: 	1194 
    -- CP-element group 1195: successors 
    -- CP-element group 1195: 	1196 
    -- CP-element group 1195: 	1197 
    -- CP-element group 1195:  members (1) 
      -- CP-element group 1195: 	 branch_block_stmt_1353/merge_stmt_2594_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1195) <= minSumDecode_CP_6680_elements(1194);
    -- CP-element group 1196:  transition  input  no-bypass 
    -- CP-element group 1196: predecessors 
    -- CP-element group 1196: 	1195 
    -- CP-element group 1196: successors 
    -- CP-element group 1196: 	1198 
    -- CP-element group 1196:  members (1) 
      -- CP-element group 1196: 	 branch_block_stmt_1353/merge_stmt_2594_PhiAck/phi_stmt_2595_ack
      -- 
    phi_stmt_2595_ack_13438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2595_ack_0, ack => minSumDecode_CP_6680_elements(1196)); -- 
    -- CP-element group 1197:  transition  input  no-bypass 
    -- CP-element group 1197: predecessors 
    -- CP-element group 1197: 	1195 
    -- CP-element group 1197: successors 
    -- CP-element group 1197: 	1198 
    -- CP-element group 1197:  members (1) 
      -- CP-element group 1197: 	 branch_block_stmt_1353/merge_stmt_2594_PhiAck/phi_stmt_2601_ack
      -- 
    phi_stmt_2601_ack_13439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2601_ack_0, ack => minSumDecode_CP_6680_elements(1197)); -- 
    -- CP-element group 1198:  join  transition  bypass 
    -- CP-element group 1198: predecessors 
    -- CP-element group 1198: 	1196 
    -- CP-element group 1198: 	1197 
    -- CP-element group 1198: successors 
    -- CP-element group 1198: 	97 
    -- CP-element group 1198:  members (1) 
      -- CP-element group 1198: 	 branch_block_stmt_1353/merge_stmt_2594_PhiAck/$exit
      -- 
    minSumDecode_cp_element_group_1198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1196) & minSumDecode_CP_6680_elements(1197);
      gj_minSumDecode_cp_element_group_1198 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1199:  transition  bypass 
    -- CP-element group 1199: predecessors 
    -- CP-element group 1199: 	818 
    -- CP-element group 1199: successors 
    -- CP-element group 1199: 	1200 
    -- CP-element group 1199:  members (2) 
      -- CP-element group 1199: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_bbx_xnphx_xi13x_xpreheader_PhiReq/$entry
      -- CP-element group 1199: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_bbx_xnphx_xi13x_xpreheader_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1199) <= minSumDecode_CP_6680_elements(818);
    -- CP-element group 1200:  place  bypass 
    -- CP-element group 1200: predecessors 
    -- CP-element group 1200: 	1199 
    -- CP-element group 1200: successors 
    -- CP-element group 1200: 	1201 
    -- CP-element group 1200:  members (1) 
      -- CP-element group 1200: 	 branch_block_stmt_1353/merge_stmt_2623_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1200) <= minSumDecode_CP_6680_elements(1199);
    -- CP-element group 1201:  transition  bypass 
    -- CP-element group 1201: predecessors 
    -- CP-element group 1201: 	1200 
    -- CP-element group 1201: successors 
    -- CP-element group 1201: 	99 
    -- CP-element group 1201:  members (3) 
      -- CP-element group 1201: 	 branch_block_stmt_1353/merge_stmt_2623_PhiAck/$entry
      -- CP-element group 1201: 	 branch_block_stmt_1353/merge_stmt_2623_PhiAck/$exit
      -- CP-element group 1201: 	 branch_block_stmt_1353/merge_stmt_2623_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1201) <= minSumDecode_CP_6680_elements(1200);
    -- CP-element group 1202:  fork  transition  output  bypass 
    -- CP-element group 1202: predecessors 
    -- CP-element group 1202: 	848 
    -- CP-element group 1202: successors 
    -- CP-element group 1202: 	1203 
    -- CP-element group 1202: 	1204 
    -- CP-element group 1202:  members (9) 
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Sample/rr
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Update/cr
      -- 
    rr_13470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1202), ack => type_cast_2629_inst_req_0); -- 
    cr_13475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1202), ack => type_cast_2629_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1202) <= minSumDecode_CP_6680_elements(848);
    -- CP-element group 1203:  transition  input  no-bypass 
    -- CP-element group 1203: predecessors 
    -- CP-element group 1203: 	1202 
    -- CP-element group 1203: successors 
    -- CP-element group 1203: 	1205 
    -- CP-element group 1203:  members (2) 
      -- CP-element group 1203: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Sample/$exit
      -- CP-element group 1203: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Sample/ra
      -- 
    ra_13471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_0, ack => minSumDecode_CP_6680_elements(1203)); -- 
    -- CP-element group 1204:  transition  input  no-bypass 
    -- CP-element group 1204: predecessors 
    -- CP-element group 1204: 	1202 
    -- CP-element group 1204: successors 
    -- CP-element group 1204: 	1205 
    -- CP-element group 1204:  members (2) 
      -- CP-element group 1204: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Update/$exit
      -- CP-element group 1204: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/Update/ca
      -- 
    ca_13476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_1, ack => minSumDecode_CP_6680_elements(1204)); -- 
    -- CP-element group 1205:  join  transition  output  bypass 
    -- CP-element group 1205: predecessors 
    -- CP-element group 1205: 	1203 
    -- CP-element group 1205: 	1204 
    -- CP-element group 1205: successors 
    -- CP-element group 1205: 	1209 
    -- CP-element group 1205:  members (6) 
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/$exit
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/$exit
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/$exit
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/$exit
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2629/SplitProtocol/$exit
      -- CP-element group 1205: 	 branch_block_stmt_1353/bbx_xnphx_xi13_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_req
      -- 
    phi_stmt_2626_req_13477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2626_req_13477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1205), ack => phi_stmt_2626_req_0); -- 
    minSumDecode_cp_element_group_1205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1203) & minSumDecode_CP_6680_elements(1204);
      gj_minSumDecode_cp_element_group_1205 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1206:  transition  bypass 
    -- CP-element group 1206: predecessors 
    -- CP-element group 1206: 	99 
    -- CP-element group 1206: successors 
    -- CP-element group 1206: 	1207 
    -- CP-element group 1206:  members (3) 
      -- CP-element group 1206: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/$entry
      -- CP-element group 1206: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/$entry
      -- CP-element group 1206: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/$entry
      -- 
    minSumDecode_CP_6680_elements(1206) <= minSumDecode_CP_6680_elements(99);
    -- CP-element group 1207:  transition  bypass 
    -- CP-element group 1207: predecessors 
    -- CP-element group 1207: 	1206 
    -- CP-element group 1207: successors 
    -- CP-element group 1207: 	1208 
    -- CP-element group 1207:  members (1) 
      -- CP-element group 1207: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/type_cast_2632_konst_delay_trans
      -- 
    -- Element group minSumDecode_CP_6680_elements(1207) is a control-delay.
    cp_element_1207_delay: control_delay_element  generic map(name => " 1207_delay", delay_value => 1)  port map(req => minSumDecode_CP_6680_elements(1206), ack => minSumDecode_CP_6680_elements(1207), clk => clk, reset =>reset);
    -- CP-element group 1208:  transition  output  bypass 
    -- CP-element group 1208: predecessors 
    -- CP-element group 1208: 	1207 
    -- CP-element group 1208: successors 
    -- CP-element group 1208: 	1209 
    -- CP-element group 1208:  members (4) 
      -- CP-element group 1208: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/$exit
      -- CP-element group 1208: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/$exit
      -- CP-element group 1208: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_sources/$exit
      -- CP-element group 1208: 	 branch_block_stmt_1353/bbx_xnphx_xi13x_xpreheader_bbx_xnphx_xi13_PhiReq/phi_stmt_2626/phi_stmt_2626_req
      -- 
    phi_stmt_2626_req_13488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2626_req_13488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1208), ack => phi_stmt_2626_req_1); -- 
    minSumDecode_CP_6680_elements(1208) <= minSumDecode_CP_6680_elements(1207);
    -- CP-element group 1209:  merge  place  bypass 
    -- CP-element group 1209: predecessors 
    -- CP-element group 1209: 	1205 
    -- CP-element group 1209: 	1208 
    -- CP-element group 1209: successors 
    -- CP-element group 1209: 	1210 
    -- CP-element group 1209:  members (1) 
      -- CP-element group 1209: 	 branch_block_stmt_1353/merge_stmt_2625_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1209) <= OrReduce(minSumDecode_CP_6680_elements(1205) & minSumDecode_CP_6680_elements(1208));
    -- CP-element group 1210:  transition  bypass 
    -- CP-element group 1210: predecessors 
    -- CP-element group 1210: 	1209 
    -- CP-element group 1210: successors 
    -- CP-element group 1210: 	1211 
    -- CP-element group 1210:  members (1) 
      -- CP-element group 1210: 	 branch_block_stmt_1353/merge_stmt_2625_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1210) <= minSumDecode_CP_6680_elements(1209);
    -- CP-element group 1211:  transition  input  no-bypass 
    -- CP-element group 1211: predecessors 
    -- CP-element group 1211: 	1210 
    -- CP-element group 1211: successors 
    -- CP-element group 1211: 	100 
    -- CP-element group 1211:  members (2) 
      -- CP-element group 1211: 	 branch_block_stmt_1353/merge_stmt_2625_PhiAck/$exit
      -- CP-element group 1211: 	 branch_block_stmt_1353/merge_stmt_2625_PhiAck/phi_stmt_2626_ack
      -- 
    phi_stmt_2626_ack_13493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2626_ack_0, ack => minSumDecode_CP_6680_elements(1211)); -- 
    -- CP-element group 1212:  transition  bypass 
    -- CP-element group 1212: predecessors 
    -- CP-element group 1212: 	849 
    -- CP-element group 1212: successors 
    -- CP-element group 1212: 	1213 
    -- CP-element group 1212:  members (2) 
      -- CP-element group 1212: 	 branch_block_stmt_1353/bbx_xnphx_xi13_send_outputx_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 1212: 	 branch_block_stmt_1353/bbx_xnphx_xi13_send_outputx_xexitx_xloopexit_PhiReq/$exit
      -- 
    minSumDecode_CP_6680_elements(1212) <= minSumDecode_CP_6680_elements(849);
    -- CP-element group 1213:  place  bypass 
    -- CP-element group 1213: predecessors 
    -- CP-element group 1213: 	1212 
    -- CP-element group 1213: successors 
    -- CP-element group 1213: 	1214 
    -- CP-element group 1213:  members (1) 
      -- CP-element group 1213: 	 branch_block_stmt_1353/merge_stmt_2683_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1213) <= minSumDecode_CP_6680_elements(1212);
    -- CP-element group 1214:  transition  bypass 
    -- CP-element group 1214: predecessors 
    -- CP-element group 1214: 	1213 
    -- CP-element group 1214: successors 
    -- CP-element group 1214: 	104 
    -- CP-element group 1214:  members (3) 
      -- CP-element group 1214: 	 branch_block_stmt_1353/merge_stmt_2683_PhiAck/$entry
      -- CP-element group 1214: 	 branch_block_stmt_1353/merge_stmt_2683_PhiAck/$exit
      -- CP-element group 1214: 	 branch_block_stmt_1353/merge_stmt_2683_PhiAck/dummy
      -- 
    minSumDecode_CP_6680_elements(1214) <= minSumDecode_CP_6680_elements(1213);
    -- CP-element group 1215:  fork  transition  output  bypass 
    -- CP-element group 1215: predecessors 
    -- CP-element group 1215: 	817 
    -- CP-element group 1215: successors 
    -- CP-element group 1215: 	1216 
    -- CP-element group 1215: 	1217 
    -- CP-element group 1215:  members (9) 
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Sample/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Sample/rr
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Update/$entry
      -- CP-element group 1215: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Update/cr
      -- 
    rr_13524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1215), ack => type_cast_2696_inst_req_0); -- 
    cr_13529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1215), ack => type_cast_2696_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1215) <= minSumDecode_CP_6680_elements(817);
    -- CP-element group 1216:  transition  input  no-bypass 
    -- CP-element group 1216: predecessors 
    -- CP-element group 1216: 	1215 
    -- CP-element group 1216: successors 
    -- CP-element group 1216: 	1218 
    -- CP-element group 1216:  members (2) 
      -- CP-element group 1216: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Sample/$exit
      -- CP-element group 1216: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Sample/ra
      -- 
    ra_13525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_0, ack => minSumDecode_CP_6680_elements(1216)); -- 
    -- CP-element group 1217:  transition  input  no-bypass 
    -- CP-element group 1217: predecessors 
    -- CP-element group 1217: 	1215 
    -- CP-element group 1217: successors 
    -- CP-element group 1217: 	1218 
    -- CP-element group 1217:  members (2) 
      -- CP-element group 1217: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Update/$exit
      -- CP-element group 1217: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/Update/ca
      -- 
    ca_13530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_1, ack => minSumDecode_CP_6680_elements(1217)); -- 
    -- CP-element group 1218:  join  transition  output  bypass 
    -- CP-element group 1218: predecessors 
    -- CP-element group 1218: 	1216 
    -- CP-element group 1218: 	1217 
    -- CP-element group 1218: successors 
    -- CP-element group 1218: 	1227 
    -- CP-element group 1218:  members (6) 
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/$exit
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/$exit
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$exit
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/$exit
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2696/SplitProtocol/$exit
      -- CP-element group 1218: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_req
      -- 
    phi_stmt_2689_req_13531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2689_req_13531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1218), ack => phi_stmt_2689_req_2); -- 
    minSumDecode_cp_element_group_1218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1216) & minSumDecode_CP_6680_elements(1217);
      gj_minSumDecode_cp_element_group_1218 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1219:  fork  transition  output  bypass 
    -- CP-element group 1219: predecessors 
    -- CP-element group 1219: 	52 
    -- CP-element group 1219: successors 
    -- CP-element group 1219: 	1220 
    -- CP-element group 1219: 	1221 
    -- CP-element group 1219:  members (9) 
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Sample/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Sample/rr
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Update/$entry
      -- CP-element group 1219: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Update/cr
      -- 
    rr_13550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1219), ack => type_cast_2694_inst_req_0); -- 
    cr_13555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1219), ack => type_cast_2694_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1219) <= minSumDecode_CP_6680_elements(52);
    -- CP-element group 1220:  transition  input  no-bypass 
    -- CP-element group 1220: predecessors 
    -- CP-element group 1220: 	1219 
    -- CP-element group 1220: successors 
    -- CP-element group 1220: 	1222 
    -- CP-element group 1220:  members (2) 
      -- CP-element group 1220: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Sample/$exit
      -- CP-element group 1220: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Sample/ra
      -- 
    ra_13551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_0, ack => minSumDecode_CP_6680_elements(1220)); -- 
    -- CP-element group 1221:  transition  input  no-bypass 
    -- CP-element group 1221: predecessors 
    -- CP-element group 1221: 	1219 
    -- CP-element group 1221: successors 
    -- CP-element group 1221: 	1222 
    -- CP-element group 1221:  members (2) 
      -- CP-element group 1221: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Update/$exit
      -- CP-element group 1221: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/Update/ca
      -- 
    ca_13556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_1, ack => minSumDecode_CP_6680_elements(1221)); -- 
    -- CP-element group 1222:  join  transition  output  bypass 
    -- CP-element group 1222: predecessors 
    -- CP-element group 1222: 	1220 
    -- CP-element group 1222: 	1221 
    -- CP-element group 1222: successors 
    -- CP-element group 1222: 	1227 
    -- CP-element group 1222:  members (6) 
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/$exit
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/$exit
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$exit
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/$exit
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2694/SplitProtocol/$exit
      -- CP-element group 1222: 	 branch_block_stmt_1353/checkIsdecodedx_xexitx_xthreadx_xthread_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_req
      -- 
    phi_stmt_2689_req_13557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2689_req_13557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1222), ack => phi_stmt_2689_req_1); -- 
    minSumDecode_cp_element_group_1222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1220) & minSumDecode_CP_6680_elements(1221);
      gj_minSumDecode_cp_element_group_1222 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1223:  fork  transition  output  bypass 
    -- CP-element group 1223: predecessors 
    -- CP-element group 1223: 	105 
    -- CP-element group 1223: successors 
    -- CP-element group 1223: 	1224 
    -- CP-element group 1223: 	1225 
    -- CP-element group 1223:  members (9) 
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Sample/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Sample/rr
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Update/$entry
      -- CP-element group 1223: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Update/cr
      -- 
    rr_13576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1223), ack => type_cast_2692_inst_req_0); -- 
    cr_13581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1223), ack => type_cast_2692_inst_req_1); -- 
    minSumDecode_CP_6680_elements(1223) <= minSumDecode_CP_6680_elements(105);
    -- CP-element group 1224:  transition  input  no-bypass 
    -- CP-element group 1224: predecessors 
    -- CP-element group 1224: 	1223 
    -- CP-element group 1224: successors 
    -- CP-element group 1224: 	1226 
    -- CP-element group 1224:  members (2) 
      -- CP-element group 1224: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Sample/$exit
      -- CP-element group 1224: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Sample/ra
      -- 
    ra_13577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_0, ack => minSumDecode_CP_6680_elements(1224)); -- 
    -- CP-element group 1225:  transition  input  no-bypass 
    -- CP-element group 1225: predecessors 
    -- CP-element group 1225: 	1223 
    -- CP-element group 1225: successors 
    -- CP-element group 1225: 	1226 
    -- CP-element group 1225:  members (2) 
      -- CP-element group 1225: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Update/$exit
      -- CP-element group 1225: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/Update/ca
      -- 
    ca_13582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_1, ack => minSumDecode_CP_6680_elements(1225)); -- 
    -- CP-element group 1226:  join  transition  output  bypass 
    -- CP-element group 1226: predecessors 
    -- CP-element group 1226: 	1224 
    -- CP-element group 1226: 	1225 
    -- CP-element group 1226: successors 
    -- CP-element group 1226: 	1227 
    -- CP-element group 1226:  members (6) 
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/$exit
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/$exit
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/$exit
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/$exit
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_sources/type_cast_2692/SplitProtocol/$exit
      -- CP-element group 1226: 	 branch_block_stmt_1353/send_outputx_xexitx_xloopexit_send_outputx_xexit_PhiReq/phi_stmt_2689/phi_stmt_2689_req
      -- 
    phi_stmt_2689_req_13583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2689_req_13583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => minSumDecode_CP_6680_elements(1226), ack => phi_stmt_2689_req_0); -- 
    minSumDecode_cp_element_group_1226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(1224) & minSumDecode_CP_6680_elements(1225);
      gj_minSumDecode_cp_element_group_1226 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1227:  merge  place  bypass 
    -- CP-element group 1227: predecessors 
    -- CP-element group 1227: 	1218 
    -- CP-element group 1227: 	1222 
    -- CP-element group 1227: 	1226 
    -- CP-element group 1227: successors 
    -- CP-element group 1227: 	1228 
    -- CP-element group 1227:  members (1) 
      -- CP-element group 1227: 	 branch_block_stmt_1353/merge_stmt_2688_PhiReqMerge
      -- 
    minSumDecode_CP_6680_elements(1227) <= OrReduce(minSumDecode_CP_6680_elements(1218) & minSumDecode_CP_6680_elements(1222) & minSumDecode_CP_6680_elements(1226));
    -- CP-element group 1228:  transition  bypass 
    -- CP-element group 1228: predecessors 
    -- CP-element group 1228: 	1227 
    -- CP-element group 1228: successors 
    -- CP-element group 1228: 	1229 
    -- CP-element group 1228:  members (1) 
      -- CP-element group 1228: 	 branch_block_stmt_1353/merge_stmt_2688_PhiAck/$entry
      -- 
    minSumDecode_CP_6680_elements(1228) <= minSumDecode_CP_6680_elements(1227);
    -- CP-element group 1229:  transition  input  no-bypass 
    -- CP-element group 1229: predecessors 
    -- CP-element group 1229: 	1228 
    -- CP-element group 1229: successors 
    -- CP-element group 1229: 	106 
    -- CP-element group 1229:  members (2) 
      -- CP-element group 1229: 	 branch_block_stmt_1353/merge_stmt_2688_PhiAck/$exit
      -- CP-element group 1229: 	 branch_block_stmt_1353/merge_stmt_2688_PhiAck/phi_stmt_2689_ack
      -- 
    phi_stmt_2689_ack_13588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2689_ack_0, ack => minSumDecode_CP_6680_elements(1229)); -- 
    -- CP-element group 1230:  transition  bypass 
    -- CP-element group 1230: predecessors 
    -- CP-element group 1230: 	2 
    -- CP-element group 1230: successors 
    -- CP-element group 1230:  members (2) 
      -- CP-element group 1230: 	 branch_block_stmt_1353/$exit
      -- CP-element group 1230: 	 $exit
      -- 
    minSumDecode_CP_6680_elements(1230) <= minSumDecode_CP_6680_elements(2);
    -- CP-element group 1231:  join  transition  bypass  pipeline-parent 
    -- CP-element group 1231: predecessors 
    -- CP-element group 1231: 	147 
    -- CP-element group 1231: 	165 
    -- CP-element group 1231: 	176 
    -- CP-element group 1231: 	181 
    -- CP-element group 1231: 	201 
    -- CP-element group 1231: successors 
    -- CP-element group 1231: 	130 
    -- CP-element group 1231:  members (2) 
      -- CP-element group 1231: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/$exit
      -- CP-element group 1231: 	 branch_block_stmt_1353/do_while_stmt_1381/do_while_stmt_1381_loop_body/phi_stmt_1383_phi_mux_ack_ps
      -- 
    minSumDecode_cp_element_group_1231: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 16,1 => 16,2 => 16,3 => 16,4 => 16);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "minSumDecode_cp_element_group_1231"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= minSumDecode_CP_6680_elements(147) & minSumDecode_CP_6680_elements(165) & minSumDecode_CP_6680_elements(176) & minSumDecode_CP_6680_elements(181) & minSumDecode_CP_6680_elements(201);
      gj_minSumDecode_cp_element_group_1231 : generic_join generic map(name => joinName, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => minSumDecode_CP_6680_elements(1231), clk => clk, reset => reset); --
    end block;
    minSumDecode_do_while_stmt_1381_terminator_7354: loop_terminator -- 
      generic map (name => " minSumDecode_do_while_stmt_1381_terminator_7354", max_iterations_in_flight =>16) 
      port map(loop_body_exit => minSumDecode_CP_6680_elements(130),loop_continue => minSumDecode_CP_6680_elements(205),loop_terminate => minSumDecode_CP_6680_elements(203),loop_back => minSumDecode_CP_6680_elements(128),loop_exit => minSumDecode_CP_6680_elements(127),clk => clk, reset => reset); -- 
    phi_stmt_1383_phi_seq_7111_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= minSumDecode_CP_6680_elements(140);
      minSumDecode_CP_6680_elements(148)<= src_sample_reqs(0);
      src_sample_acks(0)  <= minSumDecode_CP_6680_elements(152);
      minSumDecode_CP_6680_elements(149)<= src_update_reqs(0);
      src_update_acks(0)  <= minSumDecode_CP_6680_elements(153);
      minSumDecode_CP_6680_elements(141) <= phi_mux_reqs(0);
      triggers(1)  <= minSumDecode_CP_6680_elements(142);
      minSumDecode_CP_6680_elements(154)<= src_sample_reqs(1);
      src_sample_acks(1)  <= minSumDecode_CP_6680_elements(156);
      minSumDecode_CP_6680_elements(155)<= src_update_reqs(1);
      src_update_acks(1)  <= minSumDecode_CP_6680_elements(157);
      minSumDecode_CP_6680_elements(143) <= phi_mux_reqs(1);
      phi_stmt_1383_phi_seq_7111 : phi_sequencer_v2-- 
        generic map (place_capacity => 16, ntriggers => 2, name => "phi_stmt_1383_phi_seq_7111") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => minSumDecode_CP_6680_elements(135), 
          phi_sample_ack => minSumDecode_CP_6680_elements(138), 
          phi_update_req => minSumDecode_CP_6680_elements(137), 
          phi_update_ack => minSumDecode_CP_6680_elements(139), 
          phi_mux_ack => minSumDecode_CP_6680_elements(147), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_7052_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= minSumDecode_CP_6680_elements(131);
        preds(1)  <= minSumDecode_CP_6680_elements(132);
        entry_tmerge_7052 : transition_merge -- 
          generic map(name => " entry_tmerge_7052")
          port map (preds => preds, symbol_out => minSumDecode_CP_6680_elements(133));
          -- 
    end block;
    phi_stmt_1383_req_merge_7072_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= minSumDecode_CP_6680_elements(145);
        preds(1)  <= minSumDecode_CP_6680_elements(146);
        phi_stmt_1383_req_merge_7072 : transition_merge -- 
          generic map(name => " phi_stmt_1383_req_merge_7072")
          port map (preds => preds, symbol_out => minSumDecode_CP_6680_elements(144));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_Nitr_required_2685_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_Nitr_required_2685_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ebbyNo_1463_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_ebbyNo_1463_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_maxNitr_1727_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_maxNitr_1727_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncol_ind_1573_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncol_ind_1573_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncol_ind_1915_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncol_ind_1915_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_1358_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_1358_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_1422_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_1422_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_2046_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_2046_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ncols_2663_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_ncols_2663_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_nrows_2291_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_nrows_2291_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_rate_1466_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_rate_1466_word_address_0 : std_logic_vector(0 downto 0);
    signal R_iNsTr_155_2525_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_155_2525_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_155_2539_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_155_2539_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_156_2497_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_156_2497_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_160_2516_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_160_2516_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_18_1409_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_18_1409_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_33_1658_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_33_1658_scaled : std_logic_vector(9 downto 0);
    signal R_iNsTr_99_2004_resized : std_logic_vector(9 downto 0);
    signal R_iNsTr_99_2004_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi10_2635_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi10_2635_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi19_1794_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi19_1794_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi19_1799_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi19_1799_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi28_1884_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi28_1884_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi44_2118_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi44_2118_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi44_2123_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi44_2123_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi55_1970_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi55_1970_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi6_1628_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi6_1628_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi_1513_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi_1513_scaled : std_logic_vector(9 downto 0);
    signal R_indvarx_xi_1518_resized : std_logic_vector(9 downto 0);
    signal R_indvarx_xi_1518_scaled : std_logic_vector(9 downto 0);
    signal R_tmp11_2397_resized : std_logic_vector(9 downto 0);
    signal R_tmp11_2397_scaled : std_logic_vector(9 downto 0);
    signal R_tmp13_1981_resized : std_logic_vector(9 downto 0);
    signal R_tmp13_1981_scaled : std_logic_vector(9 downto 0);
    signal R_tmp4_1639_resized : std_logic_vector(9 downto 0);
    signal R_tmp4_1639_scaled : std_logic_vector(9 downto 0);
    signal R_tmp8_2383_resized : std_logic_vector(9 downto 0);
    signal R_tmp8_2383_scaled : std_logic_vector(9 downto 0);
    signal STORE_Nitr_required_2066_data_0 : std_logic_vector(15 downto 0);
    signal STORE_Nitr_required_2066_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_Nitr_required_2608_data_0 : std_logic_vector(15 downto 0);
    signal STORE_Nitr_required_2608_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_is_decoded_2041_data_0 : std_logic_vector(15 downto 0);
    signal STORE_is_decoded_2041_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_is_decoded_2169_data_0 : std_logic_vector(15 downto 0);
    signal STORE_is_decoded_2169_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_is_decoded_2224_data_0 : std_logic_vector(15 downto 0);
    signal STORE_is_decoded_2224_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_1410_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1410_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1410_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1410_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1514_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1514_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1514_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1514_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1519_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1519_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1519_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1519_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1629_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1629_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1629_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1629_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1640_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1640_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1640_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1640_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1659_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1659_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1659_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1659_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1795_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1795_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1795_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1795_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1800_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1800_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1800_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1800_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1885_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1885_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1885_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1885_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1971_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1971_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1971_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1971_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1982_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_1982_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_1982_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_1982_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2005_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2005_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2005_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2005_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2119_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2119_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2119_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2119_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2124_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2124_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2124_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2124_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2384_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2384_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2384_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2384_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2398_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2398_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2398_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2398_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2498_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2498_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2498_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2498_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2517_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2517_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2517_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2517_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2526_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2526_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2526_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2526_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2540_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2540_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2540_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2540_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2636_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_2636_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_2636_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_2636_root_address : std_logic_vector(9 downto 0);
    signal bbx_xnphx_xi_readCodeBlockx_xexit_taken_1436 : std_logic_vector(0 downto 0);
    signal colx_x02x_xi_2473 : std_logic_vector(15 downto 0);
    signal exitcond12_2031 : std_logic_vector(0 downto 0);
    signal exitcond14_1903 : std_logic_vector(0 downto 0);
    signal exitcond15_1821 : std_logic_vector(0 downto 0);
    signal exitcond16_2264 : std_logic_vector(0 downto 0);
    signal exitcond3_1680 : std_logic_vector(0 downto 0);
    signal exitcond5_2557 : std_logic_vector(0 downto 0);
    signal exitcond6_2577 : std_logic_vector(0 downto 0);
    signal exitcond_1551 : std_logic_vector(0 downto 0);
    signal iNsTr_100_2007 : std_logic_vector(31 downto 0);
    signal iNsTr_101_2011 : std_logic_vector(31 downto 0);
    signal iNsTr_102_2016 : std_logic_vector(31 downto 0);
    signal iNsTr_106_2130 : std_logic_vector(31 downto 0);
    signal iNsTr_107_2134 : std_logic_vector(63 downto 0);
    signal iNsTr_108_2140 : std_logic_vector(0 downto 0);
    signal iNsTr_111_2151 : std_logic_vector(31 downto 0);
    signal iNsTr_112_2155 : std_logic_vector(63 downto 0);
    signal iNsTr_113_2161 : std_logic_vector(0 downto 0);
    signal iNsTr_115_2195 : std_logic_vector(0 downto 0);
    signal iNsTr_11_1603 : std_logic_vector(63 downto 0);
    signal iNsTr_121_2206 : std_logic_vector(31 downto 0);
    signal iNsTr_122_2210 : std_logic_vector(63 downto 0);
    signal iNsTr_123_2216 : std_logic_vector(0 downto 0);
    signal iNsTr_130_2282 : std_logic_vector(0 downto 0);
    signal iNsTr_132_2292 : std_logic_vector(15 downto 0);
    signal iNsTr_133_2298 : std_logic_vector(0 downto 0);
    signal iNsTr_136_2309 : std_logic_vector(31 downto 0);
    signal iNsTr_137_2315 : std_logic_vector(31 downto 0);
    signal iNsTr_138_2331 : std_logic_vector(63 downto 0);
    signal iNsTr_13_1383 : std_logic_vector(7 downto 0);
    signal iNsTr_13_at_entry_1375 : std_logic_vector(7 downto 0);
    signal iNsTr_13_at_entry_1375_1387_buffered : std_logic_vector(7 downto 0);
    signal iNsTr_140_2405 : std_logic_vector(0 downto 0);
    signal iNsTr_142_2416 : std_logic_vector(15 downto 0);
    signal iNsTr_143_2421 : std_logic_vector(15 downto 0);
    signal iNsTr_145_2427 : std_logic_vector(15 downto 0);
    signal iNsTr_146_2431 : std_logic_vector(15 downto 0);
    signal iNsTr_147_2436 : std_logic_vector(15 downto 0);
    signal iNsTr_149_2439 : std_logic_vector(15 downto 0);
    signal iNsTr_14_1400 : std_logic_vector(7 downto 0);
    signal iNsTr_150_2457 : std_logic_vector(0 downto 0);
    signal iNsTr_155_2489 : std_logic_vector(63 downto 0);
    signal iNsTr_156_2495 : std_logic_vector(63 downto 0);
    signal iNsTr_157_2500 : std_logic_vector(31 downto 0);
    signal iNsTr_158_2504 : std_logic_vector(15 downto 0);
    signal iNsTr_159_2510 : std_logic_vector(15 downto 0);
    signal iNsTr_160_2514 : std_logic_vector(63 downto 0);
    signal iNsTr_161_2519 : std_logic_vector(31 downto 0);
    signal iNsTr_162_2523 : std_logic_vector(31 downto 0);
    signal iNsTr_163_2528 : std_logic_vector(31 downto 0);
    signal iNsTr_164_2532 : std_logic_vector(31 downto 0);
    signal iNsTr_165_2537 : std_logic_vector(31 downto 0);
    signal iNsTr_166_2542 : std_logic_vector(31 downto 0);
    signal iNsTr_168_2552 : std_logic_vector(15 downto 0);
    signal iNsTr_17_1403 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1407 : std_logic_vector(63 downto 0);
    signal iNsTr_19_1412 : std_logic_vector(31 downto 0);
    signal iNsTr_21_1420 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1423 : std_logic_vector(15 downto 0);
    signal iNsTr_23_1427 : std_logic_vector(31 downto 0);
    signal iNsTr_24_1432 : std_logic_vector(0 downto 0);
    signal iNsTr_26_1707 : std_logic_vector(15 downto 0);
    signal iNsTr_27_1713 : std_logic_vector(15 downto 0);
    signal iNsTr_28_1728 : std_logic_vector(15 downto 0);
    signal iNsTr_29_1733 : std_logic_vector(0 downto 0);
    signal iNsTr_2_1359 : std_logic_vector(15 downto 0);
    signal iNsTr_31_1646 : std_logic_vector(15 downto 0);
    signal iNsTr_32_1652 : std_logic_vector(15 downto 0);
    signal iNsTr_33_1656 : std_logic_vector(63 downto 0);
    signal iNsTr_34_1661 : std_logic_vector(31 downto 0);
    signal iNsTr_35_1665 : std_logic_vector(31 downto 0);
    signal iNsTr_38_1454 : std_logic_vector(0 downto 0);
    signal iNsTr_3_1365 : std_logic_vector(0 downto 0);
    signal iNsTr_40_1746 : std_logic_vector(0 downto 0);
    signal iNsTr_43_2616 : std_logic_vector(0 downto 0);
    signal iNsTr_46_1464 : std_logic_vector(31 downto 0);
    signal iNsTr_47_1467 : std_logic_vector(31 downto 0);
    signal iNsTr_48_1472 : std_logic_vector(31 downto 0);
    signal iNsTr_49_1488 : std_logic_vector(63 downto 0);
    signal iNsTr_51_1836 : std_logic_vector(0 downto 0);
    signal iNsTr_53_1769 : std_logic_vector(63 downto 0);
    signal iNsTr_55_2689 : std_logic_vector(15 downto 0);
    signal iNsTr_5_1561 : std_logic_vector(15 downto 0);
    signal iNsTr_60_1525 : std_logic_vector(31 downto 0);
    signal iNsTr_61_1531 : std_logic_vector(31 downto 0);
    signal iNsTr_62_1536 : std_logic_vector(31 downto 0);
    signal iNsTr_66_1916 : std_logic_vector(15 downto 0);
    signal iNsTr_67_1922 : std_logic_vector(0 downto 0);
    signal iNsTr_69_1859 : std_logic_vector(63 downto 0);
    signal iNsTr_6_1574 : std_logic_vector(15 downto 0);
    signal iNsTr_71_1806 : std_logic_vector(31 downto 0);
    signal iNsTr_74_2658 : std_logic_vector(31 downto 0);
    signal iNsTr_77_2664 : std_logic_vector(15 downto 0);
    signal iNsTr_78_2668 : std_logic_vector(31 downto 0);
    signal iNsTr_79_2676 : std_logic_vector(0 downto 0);
    signal iNsTr_7_1580 : std_logic_vector(0 downto 0);
    signal iNsTr_83_2047 : std_logic_vector(15 downto 0);
    signal iNsTr_84_2053 : std_logic_vector(0 downto 0);
    signal iNsTr_86_1945 : std_logic_vector(63 downto 0);
    signal iNsTr_94_2086 : std_logic_vector(63 downto 0);
    signal iNsTr_96_1988 : std_logic_vector(15 downto 0);
    signal iNsTr_97_1994 : std_logic_vector(15 downto 0);
    signal iNsTr_98_1998 : std_logic_vector(31 downto 0);
    signal iNsTr_99_2002 : std_logic_vector(63 downto 0);
    signal indvar18_1700 : std_logic_vector(15 downto 0);
    signal indvar_1725 : std_logic_vector(15 downto 0);
    signal indvarx_xi10_2626 : std_logic_vector(63 downto 0);
    signal indvarx_xi19_1785 : std_logic_vector(63 downto 0);
    signal indvarx_xi28_1875 : std_logic_vector(63 downto 0);
    signal indvarx_xi33_2369 : std_logic_vector(63 downto 0);
    signal indvarx_xi44_2109 : std_logic_vector(63 downto 0);
    signal indvarx_xi55_1961 : std_logic_vector(63 downto 0);
    signal indvarx_xi6_1619 : std_logic_vector(63 downto 0);
    signal indvarx_xi_1504 : std_logic_vector(63 downto 0);
    signal indvarx_xlcssa17_2061 : std_logic_vector(15 downto 0);
    signal indvarx_xlcssa_2595 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2592 : std_logic_vector(15 downto 0);
    signal indvarx_xnextx_xi22_1816 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi30_1898 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi38_2572 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi47_2259 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi59_2026 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi8_1675 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi_1546 : std_logic_vector(63 downto 0);
    signal ptr_deref_1414_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1414_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1414_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1414_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1414_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1414_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1524_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1524_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1524_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1524_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1524_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1538_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1538_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1538_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1538_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1538_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1538_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1645_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1645_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1645_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1645_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1645_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1664_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1664_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1664_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1664_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1664_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1667_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1667_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1667_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1667_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1667_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1667_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1805_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1805_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1805_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1805_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1805_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1808_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1808_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1808_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1808_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1808_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1808_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1889_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1889_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1889_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1889_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1889_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1889_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1987_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1987_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1987_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1987_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1987_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1997_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1997_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1997_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_1997_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_1997_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2010_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2010_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2010_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2010_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2010_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2018_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2018_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2018_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2018_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2018_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2018_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2129_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2129_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2129_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2129_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2129_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2150_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2150_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2150_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2150_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2150_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2184_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2184_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2184_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2184_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2184_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2184_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2205_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2205_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2205_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2205_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2205_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2239_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2239_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2239_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2239_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2239_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2239_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2415_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2415_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2415_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2415_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2415_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2426_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2426_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2426_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2426_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2426_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2430_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2430_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2430_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2430_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2430_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2503_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2503_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2503_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2503_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2503_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2522_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2522_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2522_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2522_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2522_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2531_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2531_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2531_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2531_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2531_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2544_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2544_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2544_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2544_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2544_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2544_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2657_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2657_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2657_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_2657_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_2657_word_offset_0 : std_logic_vector(9 downto 0);
    signal rangex_x0x_xi_2445 : std_logic_vector(15 downto 0);
    signal scevgep18x_xi_2386 : std_logic_vector(31 downto 0);
    signal scevgep5x_xi21_1802 : std_logic_vector(31 downto 0);
    signal scevgep5x_xi46_2126 : std_logic_vector(31 downto 0);
    signal scevgep5x_xi_1521 : std_logic_vector(31 downto 0);
    signal scevgep6x_xi58_1984 : std_logic_vector(31 downto 0);
    signal scevgep6x_xi_1642 : std_logic_vector(31 downto 0);
    signal scevgepx_xi11_2638 : std_logic_vector(31 downto 0);
    signal scevgepx_xi20_1797 : std_logic_vector(31 downto 0);
    signal scevgepx_xi29_1887 : std_logic_vector(31 downto 0);
    signal scevgepx_xi34_2400 : std_logic_vector(31 downto 0);
    signal scevgepx_xi45_2121 : std_logic_vector(31 downto 0);
    signal scevgepx_xi56_1973 : std_logic_vector(31 downto 0);
    signal scevgepx_xi7_1631 : std_logic_vector(31 downto 0);
    signal scevgepx_xi_1516 : std_logic_vector(31 downto 0);
    signal tmp10_2366 : std_logic_vector(63 downto 0);
    signal tmp10x_xi_2344 : std_logic_vector(63 downto 0);
    signal tmp11_2395 : std_logic_vector(63 downto 0);
    signal tmp12x_xi_2390 : std_logic_vector(31 downto 0);
    signal tmp13_1979 : std_logic_vector(63 downto 0);
    signal tmp1_2644 : std_logic_vector(63 downto 0);
    signal tmp2x_xi_2648 : std_logic_vector(31 downto 0);
    signal tmp4_1637 : std_logic_vector(63 downto 0);
    signal tmp4x_xi17_1782 : std_logic_vector(63 downto 0);
    signal tmp4x_xi26_1872 : std_logic_vector(63 downto 0);
    signal tmp4x_xi42_2099 : std_logic_vector(63 downto 0);
    signal tmp4x_xi4_1616 : std_logic_vector(63 downto 0);
    signal tmp4x_xi53_1958 : std_logic_vector(63 downto 0);
    signal tmp4x_xi_1501 : std_logic_vector(63 downto 0);
    signal tmp64_1394 : std_logic_vector(7 downto 0);
    signal tmp6x_xi_2485 : std_logic_vector(15 downto 0);
    signal tmp7_2360 : std_logic_vector(63 downto 0);
    signal tmp7x_xi_2321 : std_logic_vector(0 downto 0);
    signal tmp82_2654 : std_logic_vector(63 downto 0);
    signal tmp8_2381 : std_logic_vector(63 downto 0);
    signal tmp_2354 : std_logic_vector(63 downto 0);
    signal tmpx_xi14_1759 : std_logic_vector(0 downto 0);
    signal tmpx_xi24_1849 : std_logic_vector(0 downto 0);
    signal tmpx_xi2_1593 : std_logic_vector(0 downto 0);
    signal tmpx_xi35_2470 : std_logic_vector(15 downto 0);
    signal tmpx_xi39_2076 : std_logic_vector(0 downto 0);
    signal tmpx_xi50_1935 : std_logic_vector(0 downto 0);
    signal tmpx_xi_1478 : std_logic_vector(0 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1379_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1386_wire : std_logic_vector(7 downto 0);
    signal type_cast_1392_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1398_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1447_wire : std_logic_vector(15 downto 0);
    signal type_cast_1452_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1482_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1492_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1508_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1510_wire : std_logic_vector(63 downto 0);
    signal type_cast_1529_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1544_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1565_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1570_wire : std_logic_vector(15 downto 0);
    signal type_cast_1578_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1591_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1614_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1623_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1625_wire : std_logic_vector(63 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1650_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1673_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1693_wire : std_logic_vector(15 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1704_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1706_wire : std_logic_vector(15 downto 0);
    signal type_cast_1710_wire : std_logic_vector(15 downto 0);
    signal type_cast_1712_wire : std_logic_vector(15 downto 0);
    signal type_cast_1716_wire : std_logic_vector(15 downto 0);
    signal type_cast_1718_wire : std_logic_vector(15 downto 0);
    signal type_cast_1723_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1757_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1763_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1780_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1789_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1791_wire : std_logic_vector(63 downto 0);
    signal type_cast_1814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1834_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1847_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1853_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1863_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1870_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1879_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1881_wire : std_logic_vector(63 downto 0);
    signal type_cast_1891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1896_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1933_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1939_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1949_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1956_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1965_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1967_wire : std_logic_vector(63 downto 0);
    signal type_cast_1977_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1992_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2024_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2043_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2051_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2064_wire : std_logic_vector(15 downto 0);
    signal type_cast_2074_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2080_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2090_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2097_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2108_wire : std_logic_vector(15 downto 0);
    signal type_cast_2113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2115_wire : std_logic_vector(63 downto 0);
    signal type_cast_2138_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2159_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2171_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2179_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2181_wire : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2193_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2226_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2234_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2236_wire : std_logic_vector(15 downto 0);
    signal type_cast_2241_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2248_wire : std_logic_vector(15 downto 0);
    signal type_cast_2250_wire : std_logic_vector(15 downto 0);
    signal type_cast_2252_wire : std_logic_vector(15 downto 0);
    signal type_cast_2257_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2275_wire : std_logic_vector(15 downto 0);
    signal type_cast_2280_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2296_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2313_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2319_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2335_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2342_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2348_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2358_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2364_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2373_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2375_wire : std_logic_vector(63 downto 0);
    signal type_cast_2442_wire : std_logic_vector(15 downto 0);
    signal type_cast_2444_wire : std_logic_vector(15 downto 0);
    signal type_cast_2448_wire : std_logic_vector(15 downto 0);
    signal type_cast_2450_wire : std_logic_vector(15 downto 0);
    signal type_cast_2455_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2468_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2477_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2479_wire : std_logic_vector(15 downto 0);
    signal type_cast_2493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2508_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2550_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2570_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2590_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2598_wire : std_logic_vector(15 downto 0);
    signal type_cast_2600_wire : std_logic_vector(15 downto 0);
    signal type_cast_2604_wire : std_logic_vector(15 downto 0);
    signal type_cast_2606_wire : std_logic_vector(15 downto 0);
    signal type_cast_2614_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2629_wire : std_logic_vector(63 downto 0);
    signal type_cast_2632_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2642_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2672_wire : std_logic_vector(31 downto 0);
    signal type_cast_2674_wire : std_logic_vector(31 downto 0);
    signal type_cast_2692_wire : std_logic_vector(15 downto 0);
    signal type_cast_2694_wire : std_logic_vector(15 downto 0);
    signal type_cast_2696_wire : std_logic_vector(15 downto 0);
    signal xx_xlcssa_1444 : std_logic_vector(15 downto 0);
    signal xx_xneg1x_xi_2350 : std_logic_vector(15 downto 0);
    signal xx_xop19x_xi_2337 : std_logic_vector(63 downto 0);
    signal xx_xop5x_xi_1865 : std_logic_vector(63 downto 0);
    signal xx_xop6x_xi16_1775 : std_logic_vector(63 downto 0);
    signal xx_xop6x_xi41_2092 : std_logic_vector(63 downto 0);
    signal xx_xop6x_xi_1494 : std_logic_vector(63 downto 0);
    signal xx_xop7x_xi52_1951 : std_logic_vector(63 downto 0);
    signal xx_xop7x_xi_1609 : std_logic_vector(63 downto 0);
    signal xx_xopx_xi15_1765 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi25_1855 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi32_2327 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi3_1599 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi40_2082 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi51_1941 : std_logic_vector(15 downto 0);
    signal xx_xopx_xi_1484 : std_logic_vector(15 downto 0);
    signal xx_xph_1690 : std_logic_vector(15 downto 0);
    signal xx_xpr62_2601 : std_logic_vector(15 downto 0);
    signal xx_xpr84_2230 : std_logic_vector(15 downto 0);
    signal xx_xpr85_2102 : std_logic_vector(15 downto 0);
    signal xx_xpr87_2175 : std_logic_vector(15 downto 0);
    signal xx_xpr_2245 : std_logic_vector(15 downto 0);
    signal xx_xpre_2686 : std_logic_vector(15 downto 0);
    signal xx_xprx_xlcssa_2272 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_Nitr_required_2685_word_address_0 <= "0";
    LOAD_ebbyNo_1463_word_address_0 <= "0";
    LOAD_maxNitr_1727_word_address_0 <= "0";
    LOAD_ncol_ind_1573_word_address_0 <= "0";
    LOAD_ncol_ind_1915_word_address_0 <= "0";
    LOAD_ncols_1358_word_address_0 <= "0";
    LOAD_ncols_1422_word_address_0 <= "0";
    LOAD_ncols_2046_word_address_0 <= "0";
    LOAD_ncols_2663_word_address_0 <= "0";
    LOAD_nrows_2291_word_address_0 <= "0";
    LOAD_rate_1466_word_address_0 <= "0";
    STORE_Nitr_required_2066_word_address_0 <= "0";
    STORE_Nitr_required_2608_word_address_0 <= "0";
    STORE_is_decoded_2041_word_address_0 <= "0";
    STORE_is_decoded_2169_word_address_0 <= "0";
    STORE_is_decoded_2224_word_address_0 <= "0";
    array_obj_ref_1410_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1410_resized_base_address <= "0000000000";
    array_obj_ref_1514_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1514_resized_base_address <= "0000000000";
    array_obj_ref_1519_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1519_resized_base_address <= "0000000000";
    array_obj_ref_1629_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1629_resized_base_address <= "0000000000";
    array_obj_ref_1640_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1640_resized_base_address <= "0000000000";
    array_obj_ref_1659_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1659_resized_base_address <= "0000000000";
    array_obj_ref_1795_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1795_resized_base_address <= "0000000000";
    array_obj_ref_1800_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1800_resized_base_address <= "0000000000";
    array_obj_ref_1885_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1885_resized_base_address <= "0000000000";
    array_obj_ref_1971_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1971_resized_base_address <= "0000000000";
    array_obj_ref_1982_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_1982_resized_base_address <= "0000000000";
    array_obj_ref_2005_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2005_resized_base_address <= "0000000000";
    array_obj_ref_2119_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2119_resized_base_address <= "0000000000";
    array_obj_ref_2124_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2124_resized_base_address <= "0000000000";
    array_obj_ref_2384_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2384_resized_base_address <= "0000000000";
    array_obj_ref_2398_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2398_resized_base_address <= "0000000000";
    array_obj_ref_2498_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2498_resized_base_address <= "0000000000";
    array_obj_ref_2517_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2517_resized_base_address <= "0000000000";
    array_obj_ref_2526_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2526_resized_base_address <= "0000000000";
    array_obj_ref_2540_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2540_resized_base_address <= "0000000000";
    array_obj_ref_2636_offset_scale_factor_0 <= "0000000001";
    array_obj_ref_2636_resized_base_address <= "0000000000";
    ptr_deref_1414_word_offset_0 <= "0000000000";
    ptr_deref_1524_word_offset_0 <= "0000000000";
    ptr_deref_1538_word_offset_0 <= "0000000000";
    ptr_deref_1645_word_offset_0 <= "0000000000";
    ptr_deref_1664_word_offset_0 <= "0000000000";
    ptr_deref_1667_word_offset_0 <= "0000000000";
    ptr_deref_1805_word_offset_0 <= "0000000000";
    ptr_deref_1808_word_offset_0 <= "0000000000";
    ptr_deref_1889_word_offset_0 <= "0000000000";
    ptr_deref_1987_word_offset_0 <= "0000000000";
    ptr_deref_1997_word_offset_0 <= "0000000000";
    ptr_deref_2010_word_offset_0 <= "0000000000";
    ptr_deref_2018_word_offset_0 <= "0000000000";
    ptr_deref_2129_word_offset_0 <= "0000000000";
    ptr_deref_2150_word_offset_0 <= "0000000000";
    ptr_deref_2184_word_offset_0 <= "0000000000";
    ptr_deref_2205_word_offset_0 <= "0000000000";
    ptr_deref_2239_word_offset_0 <= "0000000000";
    ptr_deref_2415_word_offset_0 <= "0000000000";
    ptr_deref_2426_word_offset_0 <= "0000000000";
    ptr_deref_2430_word_offset_0 <= "0000000000";
    ptr_deref_2503_word_offset_0 <= "0000000000";
    ptr_deref_2522_word_offset_0 <= "0000000000";
    ptr_deref_2531_word_offset_0 <= "0000000000";
    ptr_deref_2544_word_offset_0 <= "0000000000";
    ptr_deref_2657_word_offset_0 <= "0000000000";
    type_cast_1363_wire_constant <= "0000000000000000";
    type_cast_1379_wire_constant <= "00000000";
    type_cast_1392_wire_constant <= "00000001";
    type_cast_1398_wire_constant <= "00000001";
    type_cast_1452_wire_constant <= "0000000000000000";
    type_cast_1476_wire_constant <= "0000000000000001";
    type_cast_1482_wire_constant <= "1111111111111111";
    type_cast_1492_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1508_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1529_wire_constant <= "11000000100000000000000000000000";
    type_cast_1544_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1565_wire_constant <= "0000000000000000";
    type_cast_1568_wire_constant <= "0000000000000000";
    type_cast_1578_wire_constant <= "0000000000000000";
    type_cast_1591_wire_constant <= "0000000000000001";
    type_cast_1597_wire_constant <= "1111111111111111";
    type_cast_1607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1614_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1650_wire_constant <= "1111111111111111";
    type_cast_1673_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1696_wire_constant <= "0000000000000000";
    type_cast_1704_wire_constant <= "0000000000000000";
    type_cast_1723_wire_constant <= "0000000000000001";
    type_cast_1744_wire_constant <= "0000000000000000";
    type_cast_1757_wire_constant <= "0000000000000001";
    type_cast_1763_wire_constant <= "1111111111111111";
    type_cast_1773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1780_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1789_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1834_wire_constant <= "0000000000000000";
    type_cast_1847_wire_constant <= "0000000000000001";
    type_cast_1853_wire_constant <= "1111111111111111";
    type_cast_1863_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1870_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1879_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1891_wire_constant <= "00000000000000000000000000000000";
    type_cast_1896_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1920_wire_constant <= "0000000000000000";
    type_cast_1933_wire_constant <= "0000000000000001";
    type_cast_1939_wire_constant <= "1111111111111111";
    type_cast_1949_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1956_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1965_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1977_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1992_wire_constant <= "1111111111111111";
    type_cast_2024_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2043_wire_constant <= "0000000000000001";
    type_cast_2051_wire_constant <= "0000000000000000";
    type_cast_2074_wire_constant <= "0000000000000001";
    type_cast_2080_wire_constant <= "1111111111111111";
    type_cast_2090_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2097_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2106_wire_constant <= "0000000000000001";
    type_cast_2113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2138_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2159_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2171_wire_constant <= "0000000000000000";
    type_cast_2179_wire_constant <= "0000000000000000";
    type_cast_2186_wire_constant <= "10111111100000000000000000000000";
    type_cast_2193_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2226_wire_constant <= "0000000000000000";
    type_cast_2234_wire_constant <= "0000000000000000";
    type_cast_2241_wire_constant <= "00111111100000000000000000000000";
    type_cast_2257_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2280_wire_constant <= "0000000000000001";
    type_cast_2296_wire_constant <= "0000000000000000";
    type_cast_2313_wire_constant <= "11111111111111111111111111111111";
    type_cast_2319_wire_constant <= "0000000000000001";
    type_cast_2325_wire_constant <= "1111111111111111";
    type_cast_2335_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2348_wire_constant <= "0000000000000001";
    type_cast_2358_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_2364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2455_wire_constant <= "0000000000000000";
    type_cast_2468_wire_constant <= "1111111111111111";
    type_cast_2477_wire_constant <= "0000000000000000";
    type_cast_2493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2508_wire_constant <= "1111111111111111";
    type_cast_2550_wire_constant <= "0000000000000001";
    type_cast_2570_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2590_wire_constant <= "0000000000000001";
    type_cast_2614_wire_constant <= "0000000000000000";
    type_cast_2632_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2652_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1375: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1379_wire_constant;
      req(0) <= phi_stmt_1375_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1375",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1375_ack_0,
          idata => idata,
          odata => iNsTr_13_at_entry_1375,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1375
    phi_stmt_1383: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1386_wire & iNsTr_13_at_entry_1375_1387_buffered;
      req <= phi_stmt_1383_req_0 & phi_stmt_1383_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1383",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1383_ack_0,
          idata => idata,
          odata => iNsTr_13_1383,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1383
    phi_stmt_1444: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1447_wire;
      req(0) <= phi_stmt_1444_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1444",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1444_ack_0,
          idata => idata,
          odata => xx_xlcssa_1444,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1444
    phi_stmt_1504: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1508_wire_constant & type_cast_1510_wire;
      req <= phi_stmt_1504_req_0 & phi_stmt_1504_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1504",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1504_ack_0,
          idata => idata,
          odata => indvarx_xi_1504,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1504
    phi_stmt_1561: Block -- phi operator 
      signal idata: std_logic_vector(47 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1565_wire_constant & type_cast_1568_wire_constant & type_cast_1570_wire;
      req <= phi_stmt_1561_req_0 & phi_stmt_1561_req_1 & phi_stmt_1561_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1561",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1561_ack_0,
          idata => idata,
          odata => iNsTr_5_1561,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1561
    phi_stmt_1619: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1623_wire_constant & type_cast_1625_wire;
      req <= phi_stmt_1619_req_0 & phi_stmt_1619_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1619",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1619_ack_0,
          idata => idata,
          odata => indvarx_xi6_1619,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1619
    phi_stmt_1690: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1693_wire & type_cast_1696_wire_constant;
      req <= phi_stmt_1690_req_0 & phi_stmt_1690_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1690",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1690_ack_0,
          idata => idata,
          odata => xx_xph_1690,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1690
    phi_stmt_1700: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1704_wire_constant & type_cast_1706_wire;
      req <= phi_stmt_1700_req_0 & phi_stmt_1700_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1700",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1700_ack_0,
          idata => idata,
          odata => indvar18_1700,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1700
    phi_stmt_1707: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1710_wire & type_cast_1712_wire;
      req <= phi_stmt_1707_req_0 & phi_stmt_1707_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1707",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1707_ack_0,
          idata => idata,
          odata => iNsTr_26_1707,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1707
    phi_stmt_1713: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1716_wire & type_cast_1718_wire;
      req <= phi_stmt_1713_req_0 & phi_stmt_1713_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1713",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1713_ack_0,
          idata => idata,
          odata => iNsTr_27_1713,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1713
    phi_stmt_1785: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1789_wire_constant & type_cast_1791_wire;
      req <= phi_stmt_1785_req_0 & phi_stmt_1785_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1785",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1785_ack_0,
          idata => idata,
          odata => indvarx_xi19_1785,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1785
    phi_stmt_1875: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1879_wire_constant & type_cast_1881_wire;
      req <= phi_stmt_1875_req_0 & phi_stmt_1875_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1875",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1875_ack_0,
          idata => idata,
          odata => indvarx_xi28_1875,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1875
    phi_stmt_1961: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1965_wire_constant & type_cast_1967_wire;
      req <= phi_stmt_1961_req_0 & phi_stmt_1961_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1961",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1961_ack_0,
          idata => idata,
          odata => indvarx_xi55_1961,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1961
    phi_stmt_2061: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2064_wire;
      req(0) <= phi_stmt_2061_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2061",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2061_ack_0,
          idata => idata,
          odata => indvarx_xlcssa17_2061,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2061
    phi_stmt_2102: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2106_wire_constant & type_cast_2108_wire;
      req <= phi_stmt_2102_req_0 & phi_stmt_2102_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2102",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2102_ack_0,
          idata => idata,
          odata => xx_xpr85_2102,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2102
    phi_stmt_2109: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2113_wire_constant & type_cast_2115_wire;
      req <= phi_stmt_2109_req_0 & phi_stmt_2109_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2109",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2109_ack_0,
          idata => idata,
          odata => indvarx_xi44_2109,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2109
    phi_stmt_2175: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2179_wire_constant & type_cast_2181_wire;
      req <= phi_stmt_2175_req_0 & phi_stmt_2175_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2175",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2175_ack_0,
          idata => idata,
          odata => xx_xpr87_2175,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2175
    phi_stmt_2230: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2234_wire_constant & type_cast_2236_wire;
      req <= phi_stmt_2230_req_0 & phi_stmt_2230_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2230",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2230_ack_0,
          idata => idata,
          odata => xx_xpr84_2230,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2230
    phi_stmt_2245: Block -- phi operator 
      signal idata: std_logic_vector(47 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2248_wire & type_cast_2250_wire & type_cast_2252_wire;
      req <= phi_stmt_2245_req_0 & phi_stmt_2245_req_1 & phi_stmt_2245_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2245",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2245_ack_0,
          idata => idata,
          odata => xx_xpr_2245,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2245
    phi_stmt_2272: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2275_wire;
      req(0) <= phi_stmt_2272_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2272",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2272_ack_0,
          idata => idata,
          odata => xx_xprx_xlcssa_2272,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2272
    phi_stmt_2369: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2373_wire_constant & type_cast_2375_wire;
      req <= phi_stmt_2369_req_0 & phi_stmt_2369_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2369",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2369_ack_0,
          idata => idata,
          odata => indvarx_xi33_2369,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2369
    phi_stmt_2439: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2442_wire & type_cast_2444_wire;
      req <= phi_stmt_2439_req_0 & phi_stmt_2439_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2439",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2439_ack_0,
          idata => idata,
          odata => iNsTr_149_2439,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2439
    phi_stmt_2445: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2448_wire & type_cast_2450_wire;
      req <= phi_stmt_2445_req_0 & phi_stmt_2445_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2445",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2445_ack_0,
          idata => idata,
          odata => rangex_x0x_xi_2445,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2445
    phi_stmt_2473: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2477_wire_constant & type_cast_2479_wire;
      req <= phi_stmt_2473_req_0 & phi_stmt_2473_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2473",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2473_ack_0,
          idata => idata,
          odata => colx_x02x_xi_2473,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2473
    phi_stmt_2595: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2598_wire & type_cast_2600_wire;
      req <= phi_stmt_2595_req_0 & phi_stmt_2595_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2595",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2595_ack_0,
          idata => idata,
          odata => indvarx_xlcssa_2595,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2595
    phi_stmt_2601: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2604_wire & type_cast_2606_wire;
      req <= phi_stmt_2601_req_0 & phi_stmt_2601_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2601",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2601_ack_0,
          idata => idata,
          odata => xx_xpr62_2601,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2601
    phi_stmt_2626: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2629_wire & type_cast_2632_wire_constant;
      req <= phi_stmt_2626_req_0 & phi_stmt_2626_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2626",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2626_ack_0,
          idata => idata,
          odata => indvarx_xi10_2626,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2626
    phi_stmt_2689: Block -- phi operator 
      signal idata: std_logic_vector(47 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_2692_wire & type_cast_2694_wire & type_cast_2696_wire;
      req <= phi_stmt_2689_req_0 & phi_stmt_2689_req_1 & phi_stmt_2689_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2689",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2689_ack_0,
          idata => idata,
          odata => iNsTr_55_2689,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2689
    MUX_1500_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1500_inst_req_0;
      MUX_1500_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1500_inst_req_1;
      MUX_1500_inst_ack_1<= update_ack(0);
      MUX_1500_inst: SelectSplitProtocol generic map(name => "MUX_1500_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop6x_xi_1494, y => type_cast_1499_wire_constant, sel => tmpx_xi_1478, z => tmp4x_xi_1501, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_1615_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1615_inst_req_0;
      MUX_1615_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1615_inst_req_1;
      MUX_1615_inst_ack_1<= update_ack(0);
      MUX_1615_inst: SelectSplitProtocol generic map(name => "MUX_1615_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop7x_xi_1609, y => type_cast_1614_wire_constant, sel => tmpx_xi2_1593, z => tmp4x_xi4_1616, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_1781_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1781_inst_req_0;
      MUX_1781_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1781_inst_req_1;
      MUX_1781_inst_ack_1<= update_ack(0);
      MUX_1781_inst: SelectSplitProtocol generic map(name => "MUX_1781_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop6x_xi16_1775, y => type_cast_1780_wire_constant, sel => tmpx_xi14_1759, z => tmp4x_xi17_1782, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_1871_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1871_inst_req_0;
      MUX_1871_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1871_inst_req_1;
      MUX_1871_inst_ack_1<= update_ack(0);
      MUX_1871_inst: SelectSplitProtocol generic map(name => "MUX_1871_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop5x_xi_1865, y => type_cast_1870_wire_constant, sel => tmpx_xi24_1849, z => tmp4x_xi26_1872, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_1957_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1957_inst_req_0;
      MUX_1957_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1957_inst_req_1;
      MUX_1957_inst_ack_1<= update_ack(0);
      MUX_1957_inst: SelectSplitProtocol generic map(name => "MUX_1957_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop7x_xi52_1951, y => type_cast_1956_wire_constant, sel => tmpx_xi50_1935, z => tmp4x_xi53_1958, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_2098_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_2098_inst_req_0;
      MUX_2098_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_2098_inst_req_1;
      MUX_2098_inst_ack_1<= update_ack(0);
      MUX_2098_inst: SelectSplitProtocol generic map(name => "MUX_2098_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop6x_xi41_2092, y => type_cast_2097_wire_constant, sel => tmpx_xi39_2076, z => tmp4x_xi42_2099, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    MUX_2343_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_2343_inst_req_0;
      MUX_2343_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_2343_inst_req_1;
      MUX_2343_inst_ack_1<= update_ack(0);
      MUX_2343_inst: SelectSplitProtocol generic map(name => "MUX_2343_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => xx_xop19x_xi_2337, y => type_cast_2342_wire_constant, sel => tmp7x_xi_2321, z => tmp10x_xi_2344, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    addr_of_1411_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1411_final_reg_req_0;
      addr_of_1411_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1411_final_reg_req_1;
      addr_of_1411_final_reg_ack_1<= rack(0);
      addr_of_1411_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1411_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1410_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_1412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1515_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1515_final_reg_req_0;
      addr_of_1515_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1515_final_reg_req_1;
      addr_of_1515_final_reg_ack_1<= rack(0);
      addr_of_1515_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1515_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1514_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi_1516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1520_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1520_final_reg_req_0;
      addr_of_1520_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1520_final_reg_req_1;
      addr_of_1520_final_reg_ack_1<= rack(0);
      addr_of_1520_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1520_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1519_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep5x_xi_1521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1630_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1630_final_reg_req_0;
      addr_of_1630_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1630_final_reg_req_1;
      addr_of_1630_final_reg_ack_1<= rack(0);
      addr_of_1630_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1630_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1629_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi7_1631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1641_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1641_final_reg_req_0;
      addr_of_1641_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1641_final_reg_req_1;
      addr_of_1641_final_reg_ack_1<= rack(0);
      addr_of_1641_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1641_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1640_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep6x_xi_1642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1660_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1660_final_reg_req_0;
      addr_of_1660_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1660_final_reg_req_1;
      addr_of_1660_final_reg_ack_1<= rack(0);
      addr_of_1660_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1660_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1659_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_34_1661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1796_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1796_final_reg_req_0;
      addr_of_1796_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1796_final_reg_req_1;
      addr_of_1796_final_reg_ack_1<= rack(0);
      addr_of_1796_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1796_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1795_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi20_1797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1801_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1801_final_reg_req_0;
      addr_of_1801_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1801_final_reg_req_1;
      addr_of_1801_final_reg_ack_1<= rack(0);
      addr_of_1801_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1801_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1800_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep5x_xi21_1802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1886_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1886_final_reg_req_0;
      addr_of_1886_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1886_final_reg_req_1;
      addr_of_1886_final_reg_ack_1<= rack(0);
      addr_of_1886_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1886_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1885_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi29_1887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1972_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1972_final_reg_req_0;
      addr_of_1972_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1972_final_reg_req_1;
      addr_of_1972_final_reg_ack_1<= rack(0);
      addr_of_1972_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1972_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1971_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi56_1973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1983_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1983_final_reg_req_0;
      addr_of_1983_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1983_final_reg_req_1;
      addr_of_1983_final_reg_ack_1<= rack(0);
      addr_of_1983_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1983_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1982_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep6x_xi58_1984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2006_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2006_final_reg_req_0;
      addr_of_2006_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2006_final_reg_req_1;
      addr_of_2006_final_reg_ack_1<= rack(0);
      addr_of_2006_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2006_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2005_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_100_2007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2120_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2120_final_reg_req_0;
      addr_of_2120_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2120_final_reg_req_1;
      addr_of_2120_final_reg_ack_1<= rack(0);
      addr_of_2120_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2120_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2119_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi45_2121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2125_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2125_final_reg_req_0;
      addr_of_2125_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2125_final_reg_req_1;
      addr_of_2125_final_reg_ack_1<= rack(0);
      addr_of_2125_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2125_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2124_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep5x_xi46_2126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2385_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2385_final_reg_req_0;
      addr_of_2385_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2385_final_reg_req_1;
      addr_of_2385_final_reg_ack_1<= rack(0);
      addr_of_2385_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2385_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2384_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgep18x_xi_2386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2399_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2399_final_reg_req_0;
      addr_of_2399_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2399_final_reg_req_1;
      addr_of_2399_final_reg_ack_1<= rack(0);
      addr_of_2399_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2399_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2398_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi34_2400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2499_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2499_final_reg_req_0;
      addr_of_2499_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2499_final_reg_req_1;
      addr_of_2499_final_reg_ack_1<= rack(0);
      addr_of_2499_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2499_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2498_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_157_2500,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2518_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2518_final_reg_req_0;
      addr_of_2518_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2518_final_reg_req_1;
      addr_of_2518_final_reg_ack_1<= rack(0);
      addr_of_2518_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2518_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2517_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_161_2519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2527_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2527_final_reg_req_0;
      addr_of_2527_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2527_final_reg_req_1;
      addr_of_2527_final_reg_ack_1<= rack(0);
      addr_of_2527_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2527_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2526_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_163_2528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2541_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2541_final_reg_req_0;
      addr_of_2541_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2541_final_reg_req_1;
      addr_of_2541_final_reg_ack_1<= rack(0);
      addr_of_2541_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2541_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2540_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_166_2542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2637_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2637_final_reg_req_0;
      addr_of_2637_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2637_final_reg_req_1;
      addr_of_2637_final_reg_ack_1<= rack(0);
      addr_of_2637_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2637_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2636_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => scevgepx_xi11_2638,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    iNsTr_13_at_entry_1375_1387_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= iNsTr_13_at_entry_1375_1387_buf_req_0;
      iNsTr_13_at_entry_1375_1387_buf_ack_0<= wack(0);
      rreq(0) <= iNsTr_13_at_entry_1375_1387_buf_req_1;
      iNsTr_13_at_entry_1375_1387_buf_ack_1<= rack(0);
      iNsTr_13_at_entry_1375_1387_buf : InterlockBuffer generic map ( -- 
        name => "iNsTr_13_at_entry_1375_1387_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_13_at_entry_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_13_at_entry_1375_1387_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_14_1400,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1386_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_13_1383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1419_inst_req_0;
      type_cast_1419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1419_inst_req_1;
      type_cast_1419_inst_ack_1<= rack(0);
      type_cast_1419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp64_1394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_21_1420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1426_inst_req_0;
      type_cast_1426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1426_inst_req_1;
      type_cast_1426_inst_ack_1<= rack(0);
      type_cast_1426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_22_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_23_1427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1447_inst_req_0;
      type_cast_1447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1447_inst_req_1;
      type_cast_1447_inst_ack_1<= rack(0);
      type_cast_1447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_22_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1447_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1487_inst_req_0;
      type_cast_1487_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1487_inst_req_1;
      type_cast_1487_inst_ack_1<= rack(0);
      type_cast_1487_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1487_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi_1484,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_49_1488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1510_inst_req_0;
      type_cast_1510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1510_inst_req_1;
      type_cast_1510_inst_ack_1<= rack(0);
      type_cast_1510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_1546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1510_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1570_inst_req_0;
      type_cast_1570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1570_inst_req_1;
      type_cast_1570_inst_ack_1<= rack(0);
      type_cast_1570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xlcssa_1444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1570_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1602_inst_req_0;
      type_cast_1602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1602_inst_req_1;
      type_cast_1602_inst_ack_1<= rack(0);
      type_cast_1602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi3_1599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_11_1603,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi8_1675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1625_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1655_inst_req_0;
      type_cast_1655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1655_inst_req_1;
      type_cast_1655_inst_ack_1<= rack(0);
      type_cast_1655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_32_1652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_33_1656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1693_inst_req_0;
      type_cast_1693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1693_inst_req_1;
      type_cast_1693_inst_ack_1<= rack(0);
      type_cast_1693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_6_1574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1693_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1706_inst_req_0;
      type_cast_1706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1706_inst_req_1;
      type_cast_1706_inst_ack_1<= rack(0);
      type_cast_1706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1706_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1710_inst_req_0;
      type_cast_1710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1710_inst_req_1;
      type_cast_1710_inst_ack_1<= rack(0);
      type_cast_1710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_66_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1710_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1712_inst_req_0;
      type_cast_1712_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1712_inst_req_1;
      type_cast_1712_inst_ack_1<= rack(0);
      type_cast_1712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1712_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xph_1690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1712_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1716_inst_req_0;
      type_cast_1716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1716_inst_req_1;
      type_cast_1716_inst_ack_1<= rack(0);
      type_cast_1716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_83_2047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1716_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1718_inst_req_0;
      type_cast_1718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1718_inst_req_1;
      type_cast_1718_inst_ack_1<= rack(0);
      type_cast_1718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_5_1561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1718_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1768_inst_req_0;
      type_cast_1768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1768_inst_req_1;
      type_cast_1768_inst_ack_1<= rack(0);
      type_cast_1768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi15_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_1769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1791_inst_req_0;
      type_cast_1791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1791_inst_req_1;
      type_cast_1791_inst_ack_1<= rack(0);
      type_cast_1791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi22_1816,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1791_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1858_inst_req_0;
      type_cast_1858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1858_inst_req_1;
      type_cast_1858_inst_ack_1<= rack(0);
      type_cast_1858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi25_1855,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_69_1859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1881_inst_req_0;
      type_cast_1881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1881_inst_req_1;
      type_cast_1881_inst_ack_1<= rack(0);
      type_cast_1881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi30_1898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1881_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1944_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1944_inst_req_0;
      type_cast_1944_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1944_inst_req_1;
      type_cast_1944_inst_ack_1<= rack(0);
      type_cast_1944_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1944_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi51_1941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_86_1945,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1967_inst_req_0;
      type_cast_1967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1967_inst_req_1;
      type_cast_1967_inst_ack_1<= rack(0);
      type_cast_1967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi59_2026,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1967_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2001_inst_req_0;
      type_cast_2001_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2001_inst_req_1;
      type_cast_2001_inst_ack_1<= rack(0);
      type_cast_2001_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_97_1994,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_99_2002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2064_inst_req_0;
      type_cast_2064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2064_inst_req_1;
      type_cast_2064_inst_ack_1<= rack(0);
      type_cast_2064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_1725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2064_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2085_inst_req_0;
      type_cast_2085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2085_inst_req_1;
      type_cast_2085_inst_ack_1<= rack(0);
      type_cast_2085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi40_2082,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_94_2086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2108_inst_req_0;
      type_cast_2108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2108_inst_req_1;
      type_cast_2108_inst_ack_1<= rack(0);
      type_cast_2108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr_2245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2108_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2115_inst_req_0;
      type_cast_2115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2115_inst_req_1;
      type_cast_2115_inst_ack_1<= rack(0);
      type_cast_2115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi47_2259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2181_inst_req_0;
      type_cast_2181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2181_inst_req_1;
      type_cast_2181_inst_ack_1<= rack(0);
      type_cast_2181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr85_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2181_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2236_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2236_inst_req_0;
      type_cast_2236_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2236_inst_req_1;
      type_cast_2236_inst_ack_1<= rack(0);
      type_cast_2236_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2236_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr85_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2236_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2248_inst_req_0;
      type_cast_2248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2248_inst_req_1;
      type_cast_2248_inst_ack_1<= rack(0);
      type_cast_2248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr84_2230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2248_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2250_inst_req_0;
      type_cast_2250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2250_inst_req_1;
      type_cast_2250_inst_ack_1<= rack(0);
      type_cast_2250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr85_2102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2250_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2252_inst_req_0;
      type_cast_2252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2252_inst_req_1;
      type_cast_2252_inst_ack_1<= rack(0);
      type_cast_2252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr87_2175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2252_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2275_inst_req_0;
      type_cast_2275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2275_inst_req_1;
      type_cast_2275_inst_ack_1<= rack(0);
      type_cast_2275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpr_2245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2275_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2308_inst_req_0;
      type_cast_2308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2308_inst_req_1;
      type_cast_2308_inst_ack_1<= rack(0);
      type_cast_2308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_132_2292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_136_2309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2330_inst_req_0;
      type_cast_2330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2330_inst_req_1;
      type_cast_2330_inst_ack_1<= rack(0);
      type_cast_2330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xopx_xi32_2327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_138_2331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2353_inst_req_0;
      type_cast_2353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2353_inst_req_1;
      type_cast_2353_inst_ack_1<= rack(0);
      type_cast_2353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_66_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_2354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2375_inst_req_0;
      type_cast_2375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2375_inst_req_1;
      type_cast_2375_inst_ack_1<= rack(0);
      type_cast_2375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi38_2572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2375_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2389_inst_req_0;
      type_cast_2389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2389_inst_req_1;
      type_cast_2389_inst_ack_1<= rack(0);
      type_cast_2389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xi33_2369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12x_xi_2390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2442_inst_req_0;
      type_cast_2442_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2442_inst_req_1;
      type_cast_2442_inst_ack_1<= rack(0);
      type_cast_2442_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_142_2416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2442_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2444_inst_req_0;
      type_cast_2444_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2444_inst_req_1;
      type_cast_2444_inst_ack_1<= rack(0);
      type_cast_2444_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2444_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_145_2427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2444_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2448_inst_req_0;
      type_cast_2448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2448_inst_req_1;
      type_cast_2448_inst_ack_1<= rack(0);
      type_cast_2448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_143_2421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2448_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2450_inst_req_0;
      type_cast_2450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2450_inst_req_1;
      type_cast_2450_inst_ack_1<= rack(0);
      type_cast_2450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_147_2436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2450_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2479_inst_req_0;
      type_cast_2479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2479_inst_req_1;
      type_cast_2479_inst_ack_1<= rack(0);
      type_cast_2479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_168_2552,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2479_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2488_inst_req_0;
      type_cast_2488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2488_inst_req_1;
      type_cast_2488_inst_ack_1<= rack(0);
      type_cast_2488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6x_xi_2485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_155_2489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2513_inst_req_0;
      type_cast_2513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2513_inst_req_1;
      type_cast_2513_inst_ack_1<= rack(0);
      type_cast_2513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_159_2510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_160_2514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2598_inst_req_0;
      type_cast_2598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2598_inst_req_1;
      type_cast_2598_inst_ack_1<= rack(0);
      type_cast_2598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_1725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2598_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2600_inst_req_0;
      type_cast_2600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2600_inst_req_1;
      type_cast_2600_inst_ack_1<= rack(0);
      type_cast_2600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_1725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2600_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2604_inst_req_0;
      type_cast_2604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2604_inst_req_1;
      type_cast_2604_inst_ack_1<= rack(0);
      type_cast_2604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_83_2047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2604_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2606_inst_req_0;
      type_cast_2606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2606_inst_req_1;
      type_cast_2606_inst_ack_1<= rack(0);
      type_cast_2606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_27_1713,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2629_inst_req_0;
      type_cast_2629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2629_inst_req_1;
      type_cast_2629_inst_ack_1<= rack(0);
      type_cast_2629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp82_2654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2629_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2647_inst_req_0;
      type_cast_2647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2647_inst_req_1;
      type_cast_2647_inst_ack_1<= rack(0);
      type_cast_2647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_2644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2x_xi_2648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2667_inst_req_0;
      type_cast_2667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2667_inst_req_1;
      type_cast_2667_inst_ack_1<= rack(0);
      type_cast_2667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_77_2664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_78_2668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2672_inst
    process(tmp2x_xi_2648) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := tmp2x_xi_2648(31 downto 0);
      type_cast_2672_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2674_inst
    process(iNsTr_78_2668) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := iNsTr_78_2668(31 downto 0);
      type_cast_2674_wire <= tmp_var; -- 
    end process;
    type_cast_2692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2692_inst_req_0;
      type_cast_2692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2692_inst_req_1;
      type_cast_2692_inst_ack_1<= rack(0);
      type_cast_2692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => xx_xpre_2686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2692_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2694_inst_req_0;
      type_cast_2694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2694_inst_req_1;
      type_cast_2694_inst_ack_1<= rack(0);
      type_cast_2694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xlcssa17_2061,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2694_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2696_inst_req_0;
      type_cast_2696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2696_inst_req_1;
      type_cast_2696_inst_ack_1<= rack(0);
      type_cast_2696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xlcssa_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2696_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_Nitr_required_2685_gather_scatter
    process(LOAD_Nitr_required_2685_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_Nitr_required_2685_data_0;
      ov(15 downto 0) := iv;
      xx_xpre_2686 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ebbyNo_1463_gather_scatter
    process(LOAD_ebbyNo_1463_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ebbyNo_1463_data_0;
      ov(31 downto 0) := iv;
      iNsTr_46_1464 <= ov(31 downto 0);
      --
    end process;
    -- equivalence LOAD_maxNitr_1727_gather_scatter
    process(LOAD_maxNitr_1727_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_maxNitr_1727_data_0;
      ov(15 downto 0) := iv;
      iNsTr_28_1728 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncol_ind_1573_gather_scatter
    process(LOAD_ncol_ind_1573_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncol_ind_1573_data_0;
      ov(15 downto 0) := iv;
      iNsTr_6_1574 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncol_ind_1915_gather_scatter
    process(LOAD_ncol_ind_1915_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncol_ind_1915_data_0;
      ov(15 downto 0) := iv;
      iNsTr_66_1916 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_1358_gather_scatter
    process(LOAD_ncols_1358_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_1358_data_0;
      ov(15 downto 0) := iv;
      iNsTr_2_1359 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_1422_gather_scatter
    process(LOAD_ncols_1422_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_1422_data_0;
      ov(15 downto 0) := iv;
      iNsTr_22_1423 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_2046_gather_scatter
    process(LOAD_ncols_2046_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_2046_data_0;
      ov(15 downto 0) := iv;
      iNsTr_83_2047 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_ncols_2663_gather_scatter
    process(LOAD_ncols_2663_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ncols_2663_data_0;
      ov(15 downto 0) := iv;
      iNsTr_77_2664 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_nrows_2291_gather_scatter
    process(LOAD_nrows_2291_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_nrows_2291_data_0;
      ov(15 downto 0) := iv;
      iNsTr_132_2292 <= ov(15 downto 0);
      --
    end process;
    -- equivalence LOAD_rate_1466_gather_scatter
    process(LOAD_rate_1466_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_rate_1466_data_0;
      ov(31 downto 0) := iv;
      iNsTr_47_1467 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_Nitr_required_2066_gather_scatter
    process(indvarx_xlcssa17_2061) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xlcssa17_2061;
      ov(15 downto 0) := iv;
      STORE_Nitr_required_2066_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_Nitr_required_2608_gather_scatter
    process(indvarx_xlcssa_2595) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xlcssa_2595;
      ov(15 downto 0) := iv;
      STORE_Nitr_required_2608_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_is_decoded_2041_gather_scatter
    process(type_cast_2043_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2043_wire_constant;
      ov(15 downto 0) := iv;
      STORE_is_decoded_2041_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_is_decoded_2169_gather_scatter
    process(type_cast_2171_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2171_wire_constant;
      ov(15 downto 0) := iv;
      STORE_is_decoded_2169_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence STORE_is_decoded_2224_gather_scatter
    process(type_cast_2226_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2226_wire_constant;
      ov(15 downto 0) := iv;
      STORE_is_decoded_2224_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1410_index_0_rename
    process(R_iNsTr_18_1409_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_18_1409_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_18_1409_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1410_index_0_resize
    process(iNsTr_18_1407) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_1407;
      ov := iv(9 downto 0);
      R_iNsTr_18_1409_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1410_index_offset
    process(R_iNsTr_18_1409_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_18_1409_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1410_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1410_root_address_inst
    process(array_obj_ref_1410_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1410_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1410_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1514_index_0_rename
    process(R_indvarx_xi_1513_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi_1513_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi_1513_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1514_index_0_resize
    process(indvarx_xi_1504) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi_1504;
      ov := iv(9 downto 0);
      R_indvarx_xi_1513_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1514_index_offset
    process(R_indvarx_xi_1513_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi_1513_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1514_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1514_root_address_inst
    process(array_obj_ref_1514_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1514_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1514_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_index_0_rename
    process(R_indvarx_xi_1518_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi_1518_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi_1518_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_index_0_resize
    process(indvarx_xi_1504) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi_1504;
      ov := iv(9 downto 0);
      R_indvarx_xi_1518_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_index_offset
    process(R_indvarx_xi_1518_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi_1518_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1519_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_root_address_inst
    process(array_obj_ref_1519_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1519_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1519_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_index_0_rename
    process(R_indvarx_xi6_1628_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi6_1628_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi6_1628_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_index_0_resize
    process(indvarx_xi6_1619) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi6_1619;
      ov := iv(9 downto 0);
      R_indvarx_xi6_1628_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_index_offset
    process(R_indvarx_xi6_1628_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi6_1628_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1629_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1629_root_address_inst
    process(array_obj_ref_1629_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1629_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1629_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1640_index_0_rename
    process(R_tmp4_1639_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp4_1639_resized;
      ov(9 downto 0) := iv;
      R_tmp4_1639_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1640_index_0_resize
    process(tmp4_1637) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp4_1637;
      ov := iv(9 downto 0);
      R_tmp4_1639_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1640_index_offset
    process(R_tmp4_1639_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp4_1639_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1640_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1640_root_address_inst
    process(array_obj_ref_1640_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1640_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1640_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1659_index_0_rename
    process(R_iNsTr_33_1658_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_33_1658_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_33_1658_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1659_index_0_resize
    process(iNsTr_33_1656) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_33_1656;
      ov := iv(9 downto 0);
      R_iNsTr_33_1658_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1659_index_offset
    process(R_iNsTr_33_1658_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_33_1658_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1659_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1659_root_address_inst
    process(array_obj_ref_1659_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1659_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1659_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_0_rename
    process(R_indvarx_xi19_1794_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi19_1794_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi19_1794_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_0_resize
    process(indvarx_xi19_1785) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi19_1785;
      ov := iv(9 downto 0);
      R_indvarx_xi19_1794_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_offset
    process(R_indvarx_xi19_1794_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi19_1794_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1795_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_root_address_inst
    process(array_obj_ref_1795_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1795_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1795_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1800_index_0_rename
    process(R_indvarx_xi19_1799_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi19_1799_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi19_1799_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1800_index_0_resize
    process(indvarx_xi19_1785) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi19_1785;
      ov := iv(9 downto 0);
      R_indvarx_xi19_1799_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1800_index_offset
    process(R_indvarx_xi19_1799_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi19_1799_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1800_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1800_root_address_inst
    process(array_obj_ref_1800_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1800_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1800_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1885_index_0_rename
    process(R_indvarx_xi28_1884_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi28_1884_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi28_1884_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1885_index_0_resize
    process(indvarx_xi28_1875) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi28_1875;
      ov := iv(9 downto 0);
      R_indvarx_xi28_1884_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1885_index_offset
    process(R_indvarx_xi28_1884_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi28_1884_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1885_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1885_root_address_inst
    process(array_obj_ref_1885_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1885_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1885_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1971_index_0_rename
    process(R_indvarx_xi55_1970_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi55_1970_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi55_1970_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1971_index_0_resize
    process(indvarx_xi55_1961) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi55_1961;
      ov := iv(9 downto 0);
      R_indvarx_xi55_1970_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1971_index_offset
    process(R_indvarx_xi55_1970_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi55_1970_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1971_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1971_root_address_inst
    process(array_obj_ref_1971_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1971_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1971_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_0_rename
    process(R_tmp13_1981_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp13_1981_resized;
      ov(9 downto 0) := iv;
      R_tmp13_1981_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_0_resize
    process(tmp13_1979) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp13_1979;
      ov := iv(9 downto 0);
      R_tmp13_1981_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_index_offset
    process(R_tmp13_1981_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp13_1981_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_1982_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1982_root_address_inst
    process(array_obj_ref_1982_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1982_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_1982_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2005_index_0_rename
    process(R_iNsTr_99_2004_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_99_2004_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_99_2004_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2005_index_0_resize
    process(iNsTr_99_2002) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_99_2002;
      ov := iv(9 downto 0);
      R_iNsTr_99_2004_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2005_index_offset
    process(R_iNsTr_99_2004_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_99_2004_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2005_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2005_root_address_inst
    process(array_obj_ref_2005_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2005_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2005_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2119_index_0_rename
    process(R_indvarx_xi44_2118_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi44_2118_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi44_2118_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2119_index_0_resize
    process(indvarx_xi44_2109) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi44_2109;
      ov := iv(9 downto 0);
      R_indvarx_xi44_2118_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2119_index_offset
    process(R_indvarx_xi44_2118_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi44_2118_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2119_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2119_root_address_inst
    process(array_obj_ref_2119_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2119_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2119_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2124_index_0_rename
    process(R_indvarx_xi44_2123_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi44_2123_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi44_2123_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2124_index_0_resize
    process(indvarx_xi44_2109) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi44_2109;
      ov := iv(9 downto 0);
      R_indvarx_xi44_2123_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2124_index_offset
    process(R_indvarx_xi44_2123_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi44_2123_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2124_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2124_root_address_inst
    process(array_obj_ref_2124_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2124_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2124_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2384_index_0_rename
    process(R_tmp8_2383_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp8_2383_resized;
      ov(9 downto 0) := iv;
      R_tmp8_2383_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2384_index_0_resize
    process(tmp8_2381) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp8_2381;
      ov := iv(9 downto 0);
      R_tmp8_2383_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2384_index_offset
    process(R_tmp8_2383_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp8_2383_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2384_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2384_root_address_inst
    process(array_obj_ref_2384_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2384_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2384_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2398_index_0_rename
    process(R_tmp11_2397_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp11_2397_resized;
      ov(9 downto 0) := iv;
      R_tmp11_2397_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2398_index_0_resize
    process(tmp11_2395) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp11_2395;
      ov := iv(9 downto 0);
      R_tmp11_2397_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2398_index_offset
    process(R_tmp11_2397_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp11_2397_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2398_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2398_root_address_inst
    process(array_obj_ref_2398_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2398_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2398_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2498_index_0_rename
    process(R_iNsTr_156_2497_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_156_2497_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_156_2497_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2498_index_0_resize
    process(iNsTr_156_2495) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_156_2495;
      ov := iv(9 downto 0);
      R_iNsTr_156_2497_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2498_index_offset
    process(R_iNsTr_156_2497_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_156_2497_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2498_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2498_root_address_inst
    process(array_obj_ref_2498_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2498_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2498_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2517_index_0_rename
    process(R_iNsTr_160_2516_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_160_2516_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_160_2516_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2517_index_0_resize
    process(iNsTr_160_2514) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_160_2514;
      ov := iv(9 downto 0);
      R_iNsTr_160_2516_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2517_index_offset
    process(R_iNsTr_160_2516_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_160_2516_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2517_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2517_root_address_inst
    process(array_obj_ref_2517_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2517_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2517_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2526_index_0_rename
    process(R_iNsTr_155_2525_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_155_2525_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_155_2525_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2526_index_0_resize
    process(iNsTr_155_2489) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_155_2489;
      ov := iv(9 downto 0);
      R_iNsTr_155_2525_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2526_index_offset
    process(R_iNsTr_155_2525_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_155_2525_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2526_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2526_root_address_inst
    process(array_obj_ref_2526_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2526_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2526_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2540_index_0_rename
    process(R_iNsTr_155_2539_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_155_2539_resized;
      ov(9 downto 0) := iv;
      R_iNsTr_155_2539_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2540_index_0_resize
    process(iNsTr_155_2489) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_155_2489;
      ov := iv(9 downto 0);
      R_iNsTr_155_2539_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2540_index_offset
    process(R_iNsTr_155_2539_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_iNsTr_155_2539_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2540_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2540_root_address_inst
    process(array_obj_ref_2540_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2540_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2540_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_index_0_rename
    process(R_indvarx_xi10_2635_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi10_2635_resized;
      ov(9 downto 0) := iv;
      R_indvarx_xi10_2635_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_index_0_resize
    process(indvarx_xi10_2626) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvarx_xi10_2626;
      ov := iv(9 downto 0);
      R_indvarx_xi10_2635_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_index_offset
    process(R_indvarx_xi10_2635_scaled) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvarx_xi10_2635_scaled;
      ov(9 downto 0) := iv;
      array_obj_ref_2636_final_offset <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_root_address_inst
    process(array_obj_ref_2636_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2636_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_2636_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_addr_0
    process(ptr_deref_1414_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1414_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_base_resize
    process(iNsTr_19_1412) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_1412;
      ov := iv(9 downto 0);
      ptr_deref_1414_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_gather_scatter
    process(iNsTr_17_1403) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_1403;
      ov(31 downto 0) := iv;
      ptr_deref_1414_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_root_address_inst
    process(ptr_deref_1414_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1414_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_addr_0
    process(ptr_deref_1524_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1524_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_base_resize
    process(scevgepx_xi_1516) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi_1516;
      ov := iv(9 downto 0);
      ptr_deref_1524_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_gather_scatter
    process(ptr_deref_1524_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_data_0;
      ov(31 downto 0) := iv;
      iNsTr_60_1525 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_root_address_inst
    process(ptr_deref_1524_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1524_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1538_addr_0
    process(ptr_deref_1538_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1538_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1538_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1538_base_resize
    process(scevgep5x_xi_1521) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi_1521;
      ov := iv(9 downto 0);
      ptr_deref_1538_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1538_gather_scatter
    process(iNsTr_62_1536) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_62_1536;
      ov(31 downto 0) := iv;
      ptr_deref_1538_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1538_root_address_inst
    process(ptr_deref_1538_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1538_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1538_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1645_addr_0
    process(ptr_deref_1645_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1645_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1645_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1645_base_resize
    process(scevgep6x_xi_1642) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep6x_xi_1642;
      ov := iv(9 downto 0);
      ptr_deref_1645_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1645_gather_scatter
    process(ptr_deref_1645_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1645_data_0;
      ov(15 downto 0) := iv;
      iNsTr_31_1646 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1645_root_address_inst
    process(ptr_deref_1645_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1645_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1645_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1664_addr_0
    process(ptr_deref_1664_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1664_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1664_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1664_base_resize
    process(iNsTr_34_1661) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_1661;
      ov := iv(9 downto 0);
      ptr_deref_1664_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1664_gather_scatter
    process(ptr_deref_1664_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1664_data_0;
      ov(31 downto 0) := iv;
      iNsTr_35_1665 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1664_root_address_inst
    process(ptr_deref_1664_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1664_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1664_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_addr_0
    process(ptr_deref_1667_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1667_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1667_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_base_resize
    process(scevgepx_xi7_1631) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi7_1631;
      ov := iv(9 downto 0);
      ptr_deref_1667_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_gather_scatter
    process(iNsTr_35_1665) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_1665;
      ov(31 downto 0) := iv;
      ptr_deref_1667_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1667_root_address_inst
    process(ptr_deref_1667_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1667_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1667_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1805_addr_0
    process(ptr_deref_1805_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1805_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1805_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1805_base_resize
    process(scevgepx_xi20_1797) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi20_1797;
      ov := iv(9 downto 0);
      ptr_deref_1805_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1805_gather_scatter
    process(ptr_deref_1805_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1805_data_0;
      ov(31 downto 0) := iv;
      iNsTr_71_1806 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1805_root_address_inst
    process(ptr_deref_1805_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1805_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1805_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1808_addr_0
    process(ptr_deref_1808_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1808_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1808_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1808_base_resize
    process(scevgep5x_xi21_1802) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi21_1802;
      ov := iv(9 downto 0);
      ptr_deref_1808_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1808_gather_scatter
    process(iNsTr_71_1806) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_71_1806;
      ov(31 downto 0) := iv;
      ptr_deref_1808_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1808_root_address_inst
    process(ptr_deref_1808_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1808_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1808_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_addr_0
    process(ptr_deref_1889_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1889_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1889_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_base_resize
    process(scevgepx_xi29_1887) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi29_1887;
      ov := iv(9 downto 0);
      ptr_deref_1889_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_gather_scatter
    process(type_cast_1891_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1891_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_1889_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1889_root_address_inst
    process(ptr_deref_1889_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1889_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1889_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1987_addr_0
    process(ptr_deref_1987_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1987_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1987_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1987_base_resize
    process(scevgep6x_xi58_1984) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep6x_xi58_1984;
      ov := iv(9 downto 0);
      ptr_deref_1987_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1987_gather_scatter
    process(ptr_deref_1987_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1987_data_0;
      ov(15 downto 0) := iv;
      iNsTr_96_1988 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1987_root_address_inst
    process(ptr_deref_1987_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1987_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1987_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1997_addr_0
    process(ptr_deref_1997_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1997_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_1997_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1997_base_resize
    process(scevgepx_xi56_1973) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi56_1973;
      ov := iv(9 downto 0);
      ptr_deref_1997_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1997_gather_scatter
    process(ptr_deref_1997_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1997_data_0;
      ov(31 downto 0) := iv;
      iNsTr_98_1998 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1997_root_address_inst
    process(ptr_deref_1997_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1997_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_1997_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2010_addr_0
    process(ptr_deref_2010_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2010_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2010_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2010_base_resize
    process(iNsTr_100_2007) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_100_2007;
      ov := iv(9 downto 0);
      ptr_deref_2010_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2010_gather_scatter
    process(ptr_deref_2010_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2010_data_0;
      ov(31 downto 0) := iv;
      iNsTr_101_2011 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2010_root_address_inst
    process(ptr_deref_2010_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2010_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2010_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2018_addr_0
    process(ptr_deref_2018_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2018_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2018_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2018_base_resize
    process(iNsTr_100_2007) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_100_2007;
      ov := iv(9 downto 0);
      ptr_deref_2018_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2018_gather_scatter
    process(iNsTr_102_2016) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_102_2016;
      ov(31 downto 0) := iv;
      ptr_deref_2018_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2018_root_address_inst
    process(ptr_deref_2018_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2018_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2018_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2129_addr_0
    process(ptr_deref_2129_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2129_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2129_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2129_base_resize
    process(scevgepx_xi45_2121) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi45_2121;
      ov := iv(9 downto 0);
      ptr_deref_2129_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2129_gather_scatter
    process(ptr_deref_2129_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2129_data_0;
      ov(31 downto 0) := iv;
      iNsTr_106_2130 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2129_root_address_inst
    process(ptr_deref_2129_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2129_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2129_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_addr_0
    process(ptr_deref_2150_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2150_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_base_resize
    process(scevgep5x_xi46_2126) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi46_2126;
      ov := iv(9 downto 0);
      ptr_deref_2150_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_gather_scatter
    process(ptr_deref_2150_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_data_0;
      ov(31 downto 0) := iv;
      iNsTr_111_2151 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2150_root_address_inst
    process(ptr_deref_2150_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2150_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2150_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_addr_0
    process(ptr_deref_2184_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2184_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2184_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_base_resize
    process(scevgep5x_xi46_2126) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi46_2126;
      ov := iv(9 downto 0);
      ptr_deref_2184_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_gather_scatter
    process(type_cast_2186_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2186_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_2184_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2184_root_address_inst
    process(ptr_deref_2184_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2184_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2184_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2205_addr_0
    process(ptr_deref_2205_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2205_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2205_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2205_base_resize
    process(scevgep5x_xi46_2126) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi46_2126;
      ov := iv(9 downto 0);
      ptr_deref_2205_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2205_gather_scatter
    process(ptr_deref_2205_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2205_data_0;
      ov(31 downto 0) := iv;
      iNsTr_121_2206 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2205_root_address_inst
    process(ptr_deref_2205_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2205_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2205_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2239_addr_0
    process(ptr_deref_2239_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2239_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2239_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2239_base_resize
    process(scevgep5x_xi46_2126) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep5x_xi46_2126;
      ov := iv(9 downto 0);
      ptr_deref_2239_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2239_gather_scatter
    process(type_cast_2241_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2241_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_2239_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2239_root_address_inst
    process(ptr_deref_2239_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2239_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2239_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_addr_0
    process(ptr_deref_2415_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2415_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_base_resize
    process(scevgepx_xi34_2400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi34_2400;
      ov := iv(9 downto 0);
      ptr_deref_2415_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_gather_scatter
    process(ptr_deref_2415_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_data_0;
      ov(15 downto 0) := iv;
      iNsTr_142_2416 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_root_address_inst
    process(ptr_deref_2415_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2415_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2426_addr_0
    process(ptr_deref_2426_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2426_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2426_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2426_base_resize
    process(scevgepx_xi34_2400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi34_2400;
      ov := iv(9 downto 0);
      ptr_deref_2426_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2426_gather_scatter
    process(ptr_deref_2426_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2426_data_0;
      ov(15 downto 0) := iv;
      iNsTr_145_2427 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2426_root_address_inst
    process(ptr_deref_2426_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2426_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2426_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2430_addr_0
    process(ptr_deref_2430_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2430_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2430_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2430_base_resize
    process(scevgep18x_xi_2386) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgep18x_xi_2386;
      ov := iv(9 downto 0);
      ptr_deref_2430_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2430_gather_scatter
    process(ptr_deref_2430_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2430_data_0;
      ov(15 downto 0) := iv;
      iNsTr_146_2431 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2430_root_address_inst
    process(ptr_deref_2430_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2430_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2430_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_addr_0
    process(ptr_deref_2503_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2503_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_base_resize
    process(iNsTr_157_2500) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_157_2500;
      ov := iv(9 downto 0);
      ptr_deref_2503_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_gather_scatter
    process(ptr_deref_2503_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_data_0;
      ov(15 downto 0) := iv;
      iNsTr_158_2504 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2503_root_address_inst
    process(ptr_deref_2503_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2503_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2503_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_addr_0
    process(ptr_deref_2522_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2522_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_base_resize
    process(iNsTr_161_2519) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_161_2519;
      ov := iv(9 downto 0);
      ptr_deref_2522_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_gather_scatter
    process(ptr_deref_2522_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_data_0;
      ov(31 downto 0) := iv;
      iNsTr_162_2523 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2522_root_address_inst
    process(ptr_deref_2522_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2522_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2522_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2531_addr_0
    process(ptr_deref_2531_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2531_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2531_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2531_base_resize
    process(iNsTr_163_2528) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_163_2528;
      ov := iv(9 downto 0);
      ptr_deref_2531_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2531_gather_scatter
    process(ptr_deref_2531_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2531_data_0;
      ov(31 downto 0) := iv;
      iNsTr_164_2532 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2531_root_address_inst
    process(ptr_deref_2531_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2531_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2531_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_addr_0
    process(ptr_deref_2544_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2544_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2544_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_base_resize
    process(iNsTr_166_2542) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_166_2542;
      ov := iv(9 downto 0);
      ptr_deref_2544_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_gather_scatter
    process(iNsTr_165_2537) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_165_2537;
      ov(31 downto 0) := iv;
      ptr_deref_2544_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2544_root_address_inst
    process(ptr_deref_2544_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2544_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2544_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2657_addr_0
    process(ptr_deref_2657_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2657_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_2657_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2657_base_resize
    process(scevgepx_xi11_2638) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := scevgepx_xi11_2638;
      ov := iv(9 downto 0);
      ptr_deref_2657_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2657_gather_scatter
    process(ptr_deref_2657_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2657_data_0;
      ov(31 downto 0) := iv;
      iNsTr_74_2658 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2657_root_address_inst
    process(ptr_deref_2657_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2657_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_2657_root_address <= ov(9 downto 0);
      --
    end process;
    do_while_stmt_1381_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_24_1432;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1381_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1381_branch_req_0,
          ack0 => do_while_stmt_1381_branch_ack_0,
          ack1 => do_while_stmt_1381_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1366_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_1365;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1366_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1366_branch_req_0,
          ack0 => if_stmt_1366_branch_ack_0,
          ack1 => if_stmt_1366_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1439_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= bbx_xnphx_xi_readCodeBlockx_xexit_taken_1436;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1439_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1439_branch_req_0,
          ack0 => if_stmt_1439_branch_ack_0,
          ack1 => if_stmt_1439_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1455_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_38_1454;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1455_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1455_branch_req_0,
          ack0 => if_stmt_1455_branch_ack_0,
          ack1 => if_stmt_1455_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1552_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1551;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1552_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1552_branch_req_0,
          ack0 => if_stmt_1552_branch_ack_0,
          ack1 => if_stmt_1552_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1581_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_7_1580;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1581_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1581_branch_req_0,
          ack0 => if_stmt_1581_branch_ack_0,
          ack1 => if_stmt_1581_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1681_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_1680;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1681_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1681_branch_req_0,
          ack0 => if_stmt_1681_branch_ack_0,
          ack1 => if_stmt_1681_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1734_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_29_1733;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1734_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1734_branch_req_0,
          ack0 => if_stmt_1734_branch_ack_0,
          ack1 => if_stmt_1734_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1747_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_40_1746;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1747_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1747_branch_req_0,
          ack0 => if_stmt_1747_branch_ack_0,
          ack1 => if_stmt_1747_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1822_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond15_1821;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1822_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1822_branch_req_0,
          ack0 => if_stmt_1822_branch_ack_0,
          ack1 => if_stmt_1822_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1837_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_51_1836;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1837_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1837_branch_req_0,
          ack0 => if_stmt_1837_branch_ack_0,
          ack1 => if_stmt_1837_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1904_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond14_1903;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1904_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1904_branch_req_0,
          ack0 => if_stmt_1904_branch_ack_0,
          ack1 => if_stmt_1904_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1923_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_67_1922;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1923_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1923_branch_req_0,
          ack0 => if_stmt_1923_branch_ack_0,
          ack1 => if_stmt_1923_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2032_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond12_2031;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2032_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2032_branch_req_0,
          ack0 => if_stmt_2032_branch_ack_0,
          ack1 => if_stmt_2032_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2054_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_84_2053;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2054_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2054_branch_req_0,
          ack0 => if_stmt_2054_branch_ack_0,
          ack1 => if_stmt_2054_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2141_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_108_2140;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2141_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2141_branch_req_0,
          ack0 => if_stmt_2141_branch_ack_0,
          ack1 => if_stmt_2141_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2162_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_113_2161;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2162_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2162_branch_req_0,
          ack0 => if_stmt_2162_branch_ack_0,
          ack1 => if_stmt_2162_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2196_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_115_2195;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2196_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2196_branch_req_0,
          ack0 => if_stmt_2196_branch_ack_0,
          ack1 => if_stmt_2196_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2217_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_123_2216;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2217_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2217_branch_req_0,
          ack0 => if_stmt_2217_branch_ack_0,
          ack1 => if_stmt_2217_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2265_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond16_2264;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2265_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2265_branch_req_0,
          ack0 => if_stmt_2265_branch_ack_0,
          ack1 => if_stmt_2265_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2283_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_130_2282;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2283_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2283_branch_req_0,
          ack0 => if_stmt_2283_branch_ack_0,
          ack1 => if_stmt_2283_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2299_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_133_2298;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2299_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2299_branch_req_0,
          ack0 => if_stmt_2299_branch_ack_0,
          ack1 => if_stmt_2299_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2406_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_140_2405;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2406_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2406_branch_req_0,
          ack0 => if_stmt_2406_branch_ack_0,
          ack1 => if_stmt_2406_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2458_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_150_2457;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2458_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2458_branch_req_0,
          ack0 => if_stmt_2458_branch_ack_0,
          ack1 => if_stmt_2458_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2558_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_2557;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2558_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2558_branch_req_0,
          ack0 => if_stmt_2558_branch_ack_0,
          ack1 => if_stmt_2558_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2578_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond6_2577;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2578_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2578_branch_req_0,
          ack0 => if_stmt_2578_branch_ack_0,
          ack1 => if_stmt_2578_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2617_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_43_2616;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2617_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2617_branch_req_0,
          ack0 => if_stmt_2617_branch_ack_0,
          ack1 => if_stmt_2617_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2677_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_79_2676;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2677_branch", condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2677_branch_req_0,
          ack0 => if_stmt_2677_branch_ack_0,
          ack1 => if_stmt_2677_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_f32_f32_2015_inst 
    ApFloatAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_101_2011 & iNsTr_98_1998;
      iNsTr_102_2016 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_f32_f32_2015_inst_req_0;
      ADD_f32_f32_2015_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_f32_f32_2015_inst_req_1;
      ADD_f32_f32_2015_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      ApFloatAdd_group_0_gI: SplitGuardInterface generic map(name => "ApFloatAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatAdd_group_0",
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 1,
          use_input_buffering => true,
          full_rate => false,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u16_u16_1483_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xlcssa_1444;
      xx_xopx_xi_1484 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1483_inst_req_0;
      ADD_u16_u16_1483_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1483_inst_req_1;
      ADD_u16_u16_1483_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : ADD_u16_u16_1598_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_6_1574;
      xx_xopx_xi3_1599 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1598_inst_req_0;
      ADD_u16_u16_1598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1598_inst_req_1;
      ADD_u16_u16_1598_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : ADD_u16_u16_1651_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_31_1646;
      iNsTr_32_1652 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1651_inst_req_0;
      ADD_u16_u16_1651_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1651_inst_req_1;
      ADD_u16_u16_1651_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : ADD_u16_u16_1724_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar18_1700;
      indvar_1725 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1724_inst_req_0;
      ADD_u16_u16_1724_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1724_inst_req_1;
      ADD_u16_u16_1724_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : ADD_u16_u16_1764_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_27_1713;
      xx_xopx_xi15_1765 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1764_inst_req_0;
      ADD_u16_u16_1764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1764_inst_req_1;
      ADD_u16_u16_1764_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : ADD_u16_u16_1854_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_26_1707;
      xx_xopx_xi25_1855 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1854_inst_req_0;
      ADD_u16_u16_1854_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1854_inst_req_1;
      ADD_u16_u16_1854_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ADD_u16_u16_1940_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_1916;
      xx_xopx_xi51_1941 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1940_inst_req_0;
      ADD_u16_u16_1940_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1940_inst_req_1;
      ADD_u16_u16_1940_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : ADD_u16_u16_1993_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_96_1988;
      iNsTr_97_1994 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1993_inst_req_0;
      ADD_u16_u16_1993_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1993_inst_req_1;
      ADD_u16_u16_1993_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_8_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : ADD_u16_u16_2081_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_83_2047;
      xx_xopx_xi40_2082 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2081_inst_req_0;
      ADD_u16_u16_2081_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2081_inst_req_1;
      ADD_u16_u16_2081_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_9_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : ADD_u16_u16_2326_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_132_2292;
      xx_xopx_xi32_2327 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2326_inst_req_0;
      ADD_u16_u16_2326_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2326_inst_req_1;
      ADD_u16_u16_2326_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_10_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ADD_u16_u16_2349_inst 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_1916;
      xx_xneg1x_xi_2350 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2349_inst_req_0;
      ADD_u16_u16_2349_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2349_inst_req_1;
      ADD_u16_u16_2349_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ADD_u16_u16_2469_inst 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_149_2439;
      tmpx_xi35_2470 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2469_inst_req_0;
      ADD_u16_u16_2469_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2469_inst_req_1;
      ADD_u16_u16_2469_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_12_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ADD_u16_u16_2484_inst 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmpx_xi35_2470 & colx_x02x_xi_2473;
      tmp6x_xi_2485 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2484_inst_req_0;
      ADD_u16_u16_2484_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2484_inst_req_1;
      ADD_u16_u16_2484_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ADD_u16_u16_2509_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_158_2504;
      iNsTr_159_2510 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2509_inst_req_0;
      ADD_u16_u16_2509_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2509_inst_req_1;
      ADD_u16_u16_2509_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1111111111111111",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ADD_u16_u16_2551_inst 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= colx_x02x_xi_2473;
      iNsTr_168_2552 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2551_inst_req_0;
      ADD_u16_u16_2551_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2551_inst_req_1;
      ADD_u16_u16_2551_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ADD_u16_u16_2591_inst 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar18_1700;
      indvarx_xnext_2592 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_2591_inst_req_0;
      ADD_u16_u16_2591_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_2591_inst_req_1;
      ADD_u16_u16_2591_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ADD_u32_u32_2314_inst 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_136_2309;
      iNsTr_137_2315 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2314_inst_req_0;
      ADD_u32_u32_2314_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2314_inst_req_1;
      ADD_u32_u32_2314_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ADD_u64_u64_1493_inst 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_49_1488;
      xx_xop6x_xi_1494 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1493_inst_req_0;
      ADD_u64_u64_1493_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1493_inst_req_1;
      ADD_u64_u64_1493_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_18_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ADD_u64_u64_1545_inst 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi_1504;
      indvarx_xnextx_xi_1546 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1545_inst_req_0;
      ADD_u64_u64_1545_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1545_inst_req_1;
      ADD_u64_u64_1545_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_19_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ADD_u64_u64_1608_inst 
    ApIntAdd_group_20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_11_1603;
      xx_xop7x_xi_1609 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1608_inst_req_0;
      ADD_u64_u64_1608_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1608_inst_req_1;
      ADD_u64_u64_1608_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_20_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ADD_u64_u64_1636_inst 
    ApIntAdd_group_21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi6_1619;
      tmp4_1637 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1636_inst_req_0;
      ADD_u64_u64_1636_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1636_inst_req_1;
      ADD_u64_u64_1636_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_21_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ADD_u64_u64_1674_inst 
    ApIntAdd_group_22: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi6_1619;
      indvarx_xnextx_xi8_1675 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1674_inst_req_0;
      ADD_u64_u64_1674_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1674_inst_req_1;
      ADD_u64_u64_1674_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_22_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ADD_u64_u64_1774_inst 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_53_1769;
      xx_xop6x_xi16_1775 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1774_inst_req_0;
      ADD_u64_u64_1774_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1774_inst_req_1;
      ADD_u64_u64_1774_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ADD_u64_u64_1815_inst 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi19_1785;
      indvarx_xnextx_xi22_1816 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1815_inst_req_0;
      ADD_u64_u64_1815_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1815_inst_req_1;
      ADD_u64_u64_1815_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ADD_u64_u64_1864_inst 
    ApIntAdd_group_25: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_69_1859;
      xx_xop5x_xi_1865 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1864_inst_req_0;
      ADD_u64_u64_1864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1864_inst_req_1;
      ADD_u64_u64_1864_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_25_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ADD_u64_u64_1897_inst 
    ApIntAdd_group_26: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi28_1875;
      indvarx_xnextx_xi30_1898 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1897_inst_req_0;
      ADD_u64_u64_1897_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1897_inst_req_1;
      ADD_u64_u64_1897_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_26_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ADD_u64_u64_1950_inst 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_86_1945;
      xx_xop7x_xi52_1951 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1950_inst_req_0;
      ADD_u64_u64_1950_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1950_inst_req_1;
      ADD_u64_u64_1950_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_27_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ADD_u64_u64_1978_inst 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi55_1961;
      tmp13_1979 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1978_inst_req_0;
      ADD_u64_u64_1978_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1978_inst_req_1;
      ADD_u64_u64_1978_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : ADD_u64_u64_2025_inst 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi55_1961;
      indvarx_xnextx_xi59_2026 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2025_inst_req_0;
      ADD_u64_u64_2025_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2025_inst_req_1;
      ADD_u64_u64_2025_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : ADD_u64_u64_2091_inst 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_94_2086;
      xx_xop6x_xi41_2092 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2091_inst_req_0;
      ADD_u64_u64_2091_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2091_inst_req_1;
      ADD_u64_u64_2091_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : ADD_u64_u64_2258_inst 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi44_2109;
      indvarx_xnextx_xi47_2259 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2258_inst_req_0;
      ADD_u64_u64_2258_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2258_inst_req_1;
      ADD_u64_u64_2258_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : ADD_u64_u64_2336_inst 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_138_2331;
      xx_xop19x_xi_2337 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2336_inst_req_0;
      ADD_u64_u64_2336_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2336_inst_req_1;
      ADD_u64_u64_2336_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : ADD_u64_u64_2359_inst 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp_2354;
      tmp7_2360 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2359_inst_req_0;
      ADD_u64_u64_2359_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2359_inst_req_1;
      ADD_u64_u64_2359_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000100",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : ADD_u64_u64_2365_inst 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp_2354;
      tmp10_2366 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2365_inst_req_0;
      ADD_u64_u64_2365_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2365_inst_req_1;
      ADD_u64_u64_2365_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : ADD_u64_u64_2380_inst 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp7_2360 & indvarx_xi33_2369;
      tmp8_2381 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2380_inst_req_0;
      ADD_u64_u64_2380_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2380_inst_req_1;
      ADD_u64_u64_2380_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : ADD_u64_u64_2394_inst 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp10_2366 & indvarx_xi33_2369;
      tmp11_2395 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2394_inst_req_0;
      ADD_u64_u64_2394_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2394_inst_req_1;
      ADD_u64_u64_2394_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : ADD_u64_u64_2494_inst 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_155_2489;
      iNsTr_156_2495 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2494_inst_req_0;
      ADD_u64_u64_2494_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2494_inst_req_1;
      ADD_u64_u64_2494_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000011",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : ADD_u64_u64_2571_inst 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi33_2369;
      indvarx_xnextx_xi38_2572 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2571_inst_req_0;
      ADD_u64_u64_2571_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2571_inst_req_1;
      ADD_u64_u64_2571_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : ADD_u64_u64_2643_inst 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi10_2626;
      tmp1_2644 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2643_inst_req_0;
      ADD_u64_u64_2643_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2643_inst_req_1;
      ADD_u64_u64_2643_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : ADD_u64_u64_2653_inst 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xi10_2626;
      tmp82_2654 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2653_inst_req_0;
      ADD_u64_u64_2653_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2653_inst_req_1;
      ADD_u64_u64_2653_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_40_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_40_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : ADD_u8_u8_1393_inst 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_13_1383;
      tmp64_1394 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_1393_inst_req_0;
      ADD_u8_u8_1393_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_1393_inst_req_1;
      ADD_u8_u8_1393_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : ADD_u8_u8_1399_inst 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_13_1383;
      iNsTr_14_1400 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_1399_inst_req_0;
      ADD_u8_u8_1399_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_1399_inst_req_1;
      ADD_u8_u8_1399_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : EQ_u16_u1_1364_inst 
    ApIntEq_group_43: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_2_1359;
      iNsTr_3_1365 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1364_inst_req_0;
      EQ_u16_u1_1364_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1364_inst_req_1;
      EQ_u16_u1_1364_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_43_gI: SplitGuardInterface generic map(name => "ApIntEq_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : EQ_u16_u1_1453_inst 
    ApIntEq_group_44: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xlcssa_1444;
      iNsTr_38_1454 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1453_inst_req_0;
      EQ_u16_u1_1453_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1453_inst_req_1;
      EQ_u16_u1_1453_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_44_gI: SplitGuardInterface generic map(name => "ApIntEq_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : EQ_u16_u1_1579_inst 
    ApIntEq_group_45: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_6_1574;
      iNsTr_7_1580 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1579_inst_req_0;
      EQ_u16_u1_1579_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1579_inst_req_1;
      EQ_u16_u1_1579_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_45_gI: SplitGuardInterface generic map(name => "ApIntEq_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : EQ_u16_u1_1745_inst 
    ApIntEq_group_46: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_27_1713;
      iNsTr_40_1746 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1745_inst_req_0;
      EQ_u16_u1_1745_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1745_inst_req_1;
      EQ_u16_u1_1745_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_46_gI: SplitGuardInterface generic map(name => "ApIntEq_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : EQ_u16_u1_1835_inst 
    ApIntEq_group_47: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_26_1707;
      iNsTr_51_1836 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1835_inst_req_0;
      EQ_u16_u1_1835_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1835_inst_req_1;
      EQ_u16_u1_1835_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_47_gI: SplitGuardInterface generic map(name => "ApIntEq_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : EQ_u16_u1_1921_inst 
    ApIntEq_group_48: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_1916;
      iNsTr_67_1922 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_1921_inst_req_0;
      EQ_u16_u1_1921_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_1921_inst_req_1;
      EQ_u16_u1_1921_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_48_gI: SplitGuardInterface generic map(name => "ApIntEq_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : EQ_u16_u1_2052_inst 
    ApIntEq_group_49: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_83_2047;
      iNsTr_84_2053 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2052_inst_req_0;
      EQ_u16_u1_2052_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2052_inst_req_1;
      EQ_u16_u1_2052_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_49_gI: SplitGuardInterface generic map(name => "ApIntEq_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : EQ_u16_u1_2281_inst 
    ApIntEq_group_50: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xprx_xlcssa_2272;
      iNsTr_130_2282 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2281_inst_req_0;
      EQ_u16_u1_2281_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2281_inst_req_1;
      EQ_u16_u1_2281_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_50_gI: SplitGuardInterface generic map(name => "ApIntEq_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : EQ_u16_u1_2297_inst 
    ApIntEq_group_51: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_132_2292;
      iNsTr_133_2298 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2297_inst_req_0;
      EQ_u16_u1_2297_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2297_inst_req_1;
      EQ_u16_u1_2297_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_51_gI: SplitGuardInterface generic map(name => "ApIntEq_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : EQ_u16_u1_2456_inst 
    ApIntEq_group_52: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rangex_x0x_xi_2445;
      iNsTr_150_2457 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2456_inst_req_0;
      EQ_u16_u1_2456_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2456_inst_req_1;
      EQ_u16_u1_2456_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_52_gI: SplitGuardInterface generic map(name => "ApIntEq_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : EQ_u16_u1_2556_inst 
    ApIntEq_group_53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_168_2552 & rangex_x0x_xi_2445;
      exitcond5_2557 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2556_inst_req_0;
      EQ_u16_u1_2556_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2556_inst_req_1;
      EQ_u16_u1_2556_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_53_gI: SplitGuardInterface generic map(name => "ApIntEq_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : EQ_u16_u1_2615_inst 
    ApIntEq_group_54: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xpr62_2601;
      iNsTr_43_2616 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u16_u1_2615_inst_req_0;
      EQ_u16_u1_2615_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u16_u1_2615_inst_req_1;
      EQ_u16_u1_2615_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_54_gI: SplitGuardInterface generic map(name => "ApIntEq_group_54_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : EQ_u32_u1_2404_inst 
    ApIntEq_group_55: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tmp12x_xi_2390 & iNsTr_137_2315;
      iNsTr_140_2405 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_2404_inst_req_0;
      EQ_u32_u1_2404_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_2404_inst_req_1;
      EQ_u32_u1_2404_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_55_gI: SplitGuardInterface generic map(name => "ApIntEq_group_55_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_55",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : EQ_u64_u1_1550_inst 
    ApIntEq_group_56: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi_1546 & tmp4x_xi_1501;
      exitcond_1551 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_1550_inst_req_0;
      EQ_u64_u1_1550_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_1550_inst_req_1;
      EQ_u64_u1_1550_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_56_gI: SplitGuardInterface generic map(name => "ApIntEq_group_56_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_56",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : EQ_u64_u1_1679_inst 
    ApIntEq_group_57: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi8_1675 & tmp4x_xi4_1616;
      exitcond3_1680 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_1679_inst_req_0;
      EQ_u64_u1_1679_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_1679_inst_req_1;
      EQ_u64_u1_1679_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_57_gI: SplitGuardInterface generic map(name => "ApIntEq_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : EQ_u64_u1_1820_inst 
    ApIntEq_group_58: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi22_1816 & tmp4x_xi17_1782;
      exitcond15_1821 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_1820_inst_req_0;
      EQ_u64_u1_1820_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_1820_inst_req_1;
      EQ_u64_u1_1820_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_58_gI: SplitGuardInterface generic map(name => "ApIntEq_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : EQ_u64_u1_1902_inst 
    ApIntEq_group_59: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi30_1898 & tmp4x_xi26_1872;
      exitcond14_1903 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_1902_inst_req_0;
      EQ_u64_u1_1902_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_1902_inst_req_1;
      EQ_u64_u1_1902_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_59_gI: SplitGuardInterface generic map(name => "ApIntEq_group_59_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : EQ_u64_u1_2030_inst 
    ApIntEq_group_60: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi59_2026 & tmp4x_xi53_1958;
      exitcond12_2031 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_2030_inst_req_0;
      EQ_u64_u1_2030_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_2030_inst_req_1;
      EQ_u64_u1_2030_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_60_gI: SplitGuardInterface generic map(name => "ApIntEq_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : EQ_u64_u1_2263_inst 
    ApIntEq_group_61: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi47_2259 & tmp4x_xi42_2099;
      exitcond16_2264 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_2263_inst_req_0;
      EQ_u64_u1_2263_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_2263_inst_req_1;
      EQ_u64_u1_2263_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_61_gI: SplitGuardInterface generic map(name => "ApIntEq_group_61_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : EQ_u64_u1_2576_inst 
    ApIntEq_group_62: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvarx_xnextx_xi38_2572 & tmp10x_xi_2344;
      exitcond6_2577 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u64_u1_2576_inst_req_0;
      EQ_u64_u1_2576_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u64_u1_2576_inst_req_1;
      EQ_u64_u1_2576_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_62_gI: SplitGuardInterface generic map(name => "ApIntEq_group_62_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : MUL_f32_f32_1530_inst MUL_f32_f32_1535_inst MUL_f32_f32_1471_inst 
    ApFloatMul_group_63: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_60_1525 & type_cast_1529_wire_constant & iNsTr_48_1472 & iNsTr_61_1531 & iNsTr_47_1467 & iNsTr_46_1464;
      iNsTr_61_1531 <= data_out(95 downto 64);
      iNsTr_62_1536 <= data_out(63 downto 32);
      iNsTr_48_1472 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      reqL_unguarded(2) <= MUL_f32_f32_1530_inst_req_0;
      reqL_unguarded(1) <= MUL_f32_f32_1535_inst_req_0;
      reqL_unguarded(0) <= MUL_f32_f32_1471_inst_req_0;
      MUL_f32_f32_1530_inst_ack_0 <= ackL_unguarded(2);
      MUL_f32_f32_1535_inst_ack_0 <= ackL_unguarded(1);
      MUL_f32_f32_1471_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= MUL_f32_f32_1530_inst_req_1;
      reqR_unguarded(1) <= MUL_f32_f32_1535_inst_req_1;
      reqR_unguarded(0) <= MUL_f32_f32_1471_inst_req_1;
      MUL_f32_f32_1530_inst_ack_1 <= ackR_unguarded(2);
      MUL_f32_f32_1535_inst_ack_1 <= ackR_unguarded(1);
      MUL_f32_f32_1471_inst_ack_1 <= ackR_unguarded(0);
      ApFloatMul_group_63_accessRegulator_0: access_regulator_base generic map (name => "ApFloatMul_group_63_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_63_accessRegulator_1: access_regulator_base generic map (name => "ApFloatMul_group_63_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_63_accessRegulator_2: access_regulator_base generic map (name => "ApFloatMul_group_63_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApFloatMul_group_63_gI: SplitGuardInterface generic map(name => "ApFloatMul_group_63_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatMul_group_63",
          operator_id => "ApFloatMul",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 3,
          use_input_buffering => true,
          full_rate => false,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : NOT_u1_u1_1435_inst 
    ApIntNot_group_64: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_24_1432;
      bbx_xnphx_xi_readCodeBlockx_xexit_taken_1436 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1435_inst_req_0;
      NOT_u1_u1_1435_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1435_inst_req_1;
      NOT_u1_u1_1435_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_64_gI: SplitGuardInterface generic map(name => "ApIntNot_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : SGT_f64_u1_2139_inst 
    ApFloatUgt_group_65: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_107_2134;
      iNsTr_108_2140 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2139_inst_req_0;
      SGT_f64_u1_2139_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2139_inst_req_1;
      SGT_f64_u1_2139_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUgt_group_65_gI: SplitGuardInterface generic map(name => "ApFloatUgt_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_65",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : SGT_f64_u1_2160_inst 
    ApFloatUgt_group_66: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_112_2155;
      iNsTr_113_2161 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SGT_f64_u1_2160_inst_req_0;
      SGT_f64_u1_2160_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SGT_f64_u1_2160_inst_req_1;
      SGT_f64_u1_2160_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUgt_group_66_gI: SplitGuardInterface generic map(name => "ApFloatUgt_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUgt",
          name => "ApFloatUgt_group_66",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : SLT_f64_u1_2194_inst 
    ApFloatUlt_group_67: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_107_2134;
      iNsTr_115_2195 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_2194_inst_req_0;
      SLT_f64_u1_2194_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_2194_inst_req_1;
      SLT_f64_u1_2194_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUlt_group_67_gI: SplitGuardInterface generic map(name => "ApFloatUlt_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_67",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : SLT_f64_u1_2215_inst 
    ApFloatUlt_group_68: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_122_2210;
      iNsTr_123_2216 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_f64_u1_2215_inst_req_0;
      SLT_f64_u1_2215_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_f64_u1_2215_inst_req_1;
      SLT_f64_u1_2215_inst_ack_1 <= ackR_unguarded(0);
      ApFloatUlt_group_68_gI: SplitGuardInterface generic map(name => "ApFloatUlt_group_68_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApFloatUlt",
          name => "ApFloatUlt_group_68",
          input1_is_int => false, 
          input1_characteristic_width => 11, 
          input1_mantissa_width    => 52, 
          iwidth_1  => 64,
          input2_is_int => false, 
          input2_characteristic_width => 11, 
          input2_mantissa_width => 52, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : SLT_i32_u1_2675_inst 
    ApIntSlt_group_69: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_2672_wire & type_cast_2674_wire;
      iNsTr_79_2676 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SLT_i32_u1_2675_inst_req_0;
      SLT_i32_u1_2675_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SLT_i32_u1_2675_inst_req_1;
      SLT_i32_u1_2675_inst_ack_1 <= ackR_unguarded(0);
      ApIntSlt_group_69_gI: SplitGuardInterface generic map(name => "ApIntSlt_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          name => "ApIntSlt_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : SUB_f32_f32_2536_inst 
    ApFloatSub_group_70: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_162_2523 & iNsTr_164_2532;
      iNsTr_165_2537 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_f32_f32_2536_inst_req_0;
      SUB_f32_f32_2536_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_f32_f32_2536_inst_req_1;
      SUB_f32_f32_2536_inst_ack_1 <= ackR_unguarded(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      ApFloatSub_group_70_gI: SplitGuardInterface generic map(name => "ApFloatSub_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          name => "ApFloatSub_group_70",
          operator_id => "ApFloatSub",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 1,
          use_input_buffering => true,
          full_rate => false,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : SUB_u16_u16_2420_inst 
    ApIntSub_group_71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xneg1x_xi_2350 & iNsTr_142_2416;
      iNsTr_143_2421 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2420_inst_req_0;
      SUB_u16_u16_2420_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2420_inst_req_1;
      SUB_u16_u16_2420_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_71_gI: SplitGuardInterface generic map(name => "ApIntSub_group_71_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : SUB_u16_u16_2435_inst 
    ApIntSub_group_72: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_146_2431 & iNsTr_145_2427;
      iNsTr_147_2436 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2435_inst_req_0;
      SUB_u16_u16_2435_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2435_inst_req_1;
      SUB_u16_u16_2435_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_72_gI: SplitGuardInterface generic map(name => "ApIntSub_group_72_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : UGT_u16_u1_1477_inst 
    ApIntUgt_group_73: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= xx_xlcssa_1444;
      tmpx_xi_1478 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_1477_inst_req_0;
      UGT_u16_u1_1477_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_1477_inst_req_1;
      UGT_u16_u1_1477_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_73_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_73_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : UGT_u16_u1_1592_inst 
    ApIntUgt_group_74: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_6_1574;
      tmpx_xi2_1593 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_1592_inst_req_0;
      UGT_u16_u1_1592_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_1592_inst_req_1;
      UGT_u16_u1_1592_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_74_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_74_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_74",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : UGT_u16_u1_1758_inst 
    ApIntUgt_group_75: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_27_1713;
      tmpx_xi14_1759 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_1758_inst_req_0;
      UGT_u16_u1_1758_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_1758_inst_req_1;
      UGT_u16_u1_1758_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_75_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_75_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_75",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : UGT_u16_u1_1848_inst 
    ApIntUgt_group_76: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_26_1707;
      tmpx_xi24_1849 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_1848_inst_req_0;
      UGT_u16_u1_1848_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_1848_inst_req_1;
      UGT_u16_u1_1848_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_76_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_76_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_76",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : UGT_u16_u1_1934_inst 
    ApIntUgt_group_77: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_66_1916;
      tmpx_xi50_1935 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_1934_inst_req_0;
      UGT_u16_u1_1934_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_1934_inst_req_1;
      UGT_u16_u1_1934_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_77_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_77_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_77",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : UGT_u16_u1_2075_inst 
    ApIntUgt_group_78: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_83_2047;
      tmpx_xi39_2076 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_2075_inst_req_0;
      UGT_u16_u1_2075_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_2075_inst_req_1;
      UGT_u16_u1_2075_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_78_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_78_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_78",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : UGT_u16_u1_2320_inst 
    ApIntUgt_group_79: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_132_2292;
      tmp7x_xi_2321 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= UGT_u16_u1_2320_inst_req_0;
      UGT_u16_u1_2320_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= UGT_u16_u1_2320_inst_req_1;
      UGT_u16_u1_2320_inst_ack_1 <= ackR_unguarded(0);
      ApIntUgt_group_79_gI: SplitGuardInterface generic map(name => "ApIntUgt_group_79_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          name => "ApIntUgt_group_79",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : ULT_u16_u1_1732_inst 
    ApIntUlt_group_80: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= indvar_1725 & iNsTr_28_1728;
      iNsTr_29_1733 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u16_u1_1732_inst_req_0;
      ULT_u16_u1_1732_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u16_u1_1732_inst_req_1;
      ULT_u16_u1_1732_inst_ack_1 <= ackR_unguarded(0);
      ApIntUlt_group_80_gI: SplitGuardInterface generic map(name => "ApIntUlt_group_80_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_80",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : ULT_u32_u1_1431_inst 
    ApIntUlt_group_81: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_21_1420 & iNsTr_23_1427;
      iNsTr_24_1432 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ULT_u32_u1_1431_inst_req_0;
      ULT_u32_u1_1431_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ULT_u32_u1_1431_inst_req_1;
      ULT_u32_u1_1431_inst_ack_1 <= ackR_unguarded(0);
      ApIntUlt_group_81_gI: SplitGuardInterface generic map(name => "ApIntUlt_group_81_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          name => "ApIntUlt_group_81",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : type_cast_2133_inst 
    ApFloatResize_group_82: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_106_2130;
      iNsTr_107_2134 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2133_inst_req_0;
      type_cast_2133_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2133_inst_req_1;
      type_cast_2133_inst_ack_1 <= ackR_unguarded(0);
      ApFloatResize_group_82_gI: SplitGuardInterface generic map(name => "ApFloatResize_group_82_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApFloatResize_group_82",
          operator_id => "ApFloatResize",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 1,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : type_cast_2154_inst 
    ApFloatResize_group_83: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_111_2151;
      iNsTr_112_2155 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2154_inst_req_0;
      type_cast_2154_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2154_inst_req_1;
      type_cast_2154_inst_ack_1 <= ackR_unguarded(0);
      ApFloatResize_group_83_gI: SplitGuardInterface generic map(name => "ApFloatResize_group_83_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApFloatResize_group_83",
          operator_id => "ApFloatResize",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 1,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : type_cast_2209_inst 
    ApFloatResize_group_84: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= iNsTr_121_2206;
      iNsTr_122_2210 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= type_cast_2209_inst_req_0;
      type_cast_2209_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= type_cast_2209_inst_req_1;
      type_cast_2209_inst_ack_1 <= ackR_unguarded(0);
      ApFloatResize_group_84_gI: SplitGuardInterface generic map(name => "ApFloatResize_group_84_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApFloatResize_group_84",
          operator_id => "ApFloatResize",
          input1_is_int => false, 
          input1_characteristic_width => 8, 
          input1_mantissa_width    => 23, 
          iwidth_1  => 32,
          input2_is_int => false, 
          input2_characteristic_width => 8, 
          input2_mantissa_width => 23, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => false,
          output_characteristic_width  => 11, 
          output_mantissa_width => 52, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 1,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared load operator group (0) : LOAD_Nitr_required_2685_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_Nitr_required_2685_load_0_req_0;
      LOAD_Nitr_required_2685_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_Nitr_required_2685_load_0_req_1;
      LOAD_Nitr_required_2685_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_Nitr_required_2685_word_address_0;
      LOAD_Nitr_required_2685_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_ebbyNo_1463_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_ebbyNo_1463_load_0_req_0;
      LOAD_ebbyNo_1463_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ebbyNo_1463_load_0_req_1;
      LOAD_ebbyNo_1463_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ebbyNo_1463_word_address_0;
      LOAD_ebbyNo_1463_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_maxNitr_1727_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_maxNitr_1727_load_0_req_0;
      LOAD_maxNitr_1727_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_maxNitr_1727_load_0_req_1;
      LOAD_maxNitr_1727_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_maxNitr_1727_word_address_0;
      LOAD_maxNitr_1727_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : LOAD_ncol_ind_1915_load_0 LOAD_ncol_ind_1573_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= LOAD_ncol_ind_1915_load_0_req_0;
      reqL_unguarded(0) <= LOAD_ncol_ind_1573_load_0_req_0;
      LOAD_ncol_ind_1915_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_ncol_ind_1573_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_ncol_ind_1915_load_0_req_1;
      reqR_unguarded(0) <= LOAD_ncol_ind_1573_load_0_req_1;
      LOAD_ncol_ind_1915_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_ncol_ind_1573_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncol_ind_1915_word_address_0 & LOAD_ncol_ind_1573_word_address_0;
      LOAD_ncol_ind_1915_data_0 <= data_out(31 downto 16);
      LOAD_ncol_ind_1573_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(15 downto 0),
          mtag => memory_space_10_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : LOAD_ncols_1358_load_0 LOAD_ncols_2046_load_0 LOAD_ncols_1422_load_0 LOAD_ncols_2663_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 2, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 4, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= LOAD_ncols_1358_load_0_req_0;
      reqL_unguarded(2) <= LOAD_ncols_2046_load_0_req_0;
      reqL_unguarded(1) <= LOAD_ncols_1422_load_0_req_0;
      reqL_unguarded(0) <= LOAD_ncols_2663_load_0_req_0;
      LOAD_ncols_1358_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_ncols_2046_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_ncols_1422_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_ncols_2663_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= LOAD_ncols_1358_load_0_req_1;
      reqR_unguarded(2) <= LOAD_ncols_2046_load_0_req_1;
      reqR_unguarded(1) <= LOAD_ncols_1422_load_0_req_1;
      reqR_unguarded(0) <= LOAD_ncols_2663_load_0_req_1;
      LOAD_ncols_1358_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_ncols_2046_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_ncols_1422_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_ncols_2663_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ncols_1358_word_address_0 & LOAD_ncols_2046_word_address_0 & LOAD_ncols_1422_word_address_0 & LOAD_ncols_2663_word_address_0;
      LOAD_ncols_1358_data_0 <= data_out(63 downto 48);
      LOAD_ncols_2046_data_0 <= data_out(47 downto 32);
      LOAD_ncols_1422_data_0 <= data_out(31 downto 16);
      LOAD_ncols_2663_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 1,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(0),
          mack => memory_space_11_lr_ack(0),
          maddr => memory_space_11_lr_addr(0 downto 0),
          mtag => memory_space_11_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(0),
          mack => memory_space_11_lc_ack(0),
          mdata => memory_space_11_lc_data(15 downto 0),
          mtag => memory_space_11_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : LOAD_nrows_2291_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_nrows_2291_load_0_req_0;
      LOAD_nrows_2291_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_nrows_2291_load_0_req_1;
      LOAD_nrows_2291_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_nrows_2291_word_address_0;
      LOAD_nrows_2291_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_12_lr_req(0),
          mack => memory_space_12_lr_ack(0),
          maddr => memory_space_12_lr_addr(0 downto 0),
          mtag => memory_space_12_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_12_lc_req(0),
          mack => memory_space_12_lc_ack(0),
          mdata => memory_space_12_lc_data(15 downto 0),
          mtag => memory_space_12_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : LOAD_rate_1466_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_rate_1466_load_0_req_0;
      LOAD_rate_1466_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_rate_1466_load_0_req_1;
      LOAD_rate_1466_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_rate_1466_word_address_0;
      LOAD_rate_1466_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_13_lr_req(0),
          mack => memory_space_13_lr_ack(0),
          maddr => memory_space_13_lr_addr(0 downto 0),
          mtag => memory_space_13_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_13_lc_req(0),
          mack => memory_space_13_lc_ack(0),
          mdata => memory_space_13_lc_data(31 downto 0),
          mtag => memory_space_13_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_2205_load_0 ptr_deref_1524_load_0 ptr_deref_2150_load_0 ptr_deref_2657_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_2205_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1524_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2150_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2657_load_0_req_0;
      ptr_deref_2205_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1524_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2150_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2657_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_2205_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1524_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2150_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2657_load_0_req_1;
      ptr_deref_2205_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1524_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2150_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2657_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup7_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup7_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup7_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup7_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup7_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup7_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup7_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup7_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup7_gI: SplitGuardInterface generic map(name => "LoadGroup7_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2205_word_address_0 & ptr_deref_1524_word_address_0 & ptr_deref_2150_word_address_0 & ptr_deref_2657_word_address_0;
      ptr_deref_2205_data_0 <= data_out(127 downto 96);
      ptr_deref_1524_data_0 <= data_out(95 downto 64);
      ptr_deref_2150_data_0 <= data_out(63 downto 32);
      ptr_deref_2657_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup7", addr_width => 10,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(9 downto 0),
          mtag => memory_space_3_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup7 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : ptr_deref_1987_load_0 ptr_deref_1645_load_0 ptr_deref_2415_load_0 ptr_deref_2426_load_0 ptr_deref_2430_load_0 ptr_deref_2503_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(59 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_1987_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1645_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2415_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_2426_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2430_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2503_load_0_req_0;
      ptr_deref_1987_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1645_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2415_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_2426_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2430_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2503_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_1987_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1645_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2415_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_2426_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2430_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2503_load_0_req_1;
      ptr_deref_1987_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1645_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2415_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_2426_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2430_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2503_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup8_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup8_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup8_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup8_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup8_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup8_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup8_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup8_gI: SplitGuardInterface generic map(name => "LoadGroup8_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1987_word_address_0 & ptr_deref_1645_word_address_0 & ptr_deref_2415_word_address_0 & ptr_deref_2426_word_address_0 & ptr_deref_2430_word_address_0 & ptr_deref_2503_word_address_0;
      ptr_deref_1987_data_0 <= data_out(95 downto 80);
      ptr_deref_1645_data_0 <= data_out(79 downto 64);
      ptr_deref_2415_data_0 <= data_out(63 downto 48);
      ptr_deref_2426_data_0 <= data_out(47 downto 32);
      ptr_deref_2430_data_0 <= data_out(31 downto 16);
      ptr_deref_2503_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup8", addr_width => 10,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 4,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(9 downto 0),
          mtag => memory_space_8_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup8 load-complete ",
        data_width => 16,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : ptr_deref_1664_load_0 ptr_deref_1805_load_0 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(19 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1664_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1805_load_0_req_0;
      ptr_deref_1664_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1805_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1664_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1805_load_0_req_1;
      ptr_deref_1664_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1805_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup9_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup9_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup9_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup9_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup9_gI: SplitGuardInterface generic map(name => "LoadGroup9_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1664_word_address_0 & ptr_deref_1805_word_address_0;
      ptr_deref_1664_data_0 <= data_out(63 downto 32);
      ptr_deref_1805_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup9", addr_width => 10,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(9 downto 0),
          mtag => memory_space_2_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup9 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared load operator group (10) : ptr_deref_2531_load_0 ptr_deref_1997_load_0 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(19 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2531_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1997_load_0_req_0;
      ptr_deref_2531_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1997_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2531_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1997_load_0_req_1;
      ptr_deref_2531_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1997_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup10_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup10_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup10_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup10_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup10_gI: SplitGuardInterface generic map(name => "LoadGroup10_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2531_word_address_0 & ptr_deref_1997_word_address_0;
      ptr_deref_2531_data_0 <= data_out(63 downto 32);
      ptr_deref_1997_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup10", addr_width => 10,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(9 downto 0),
          mtag => memory_space_5_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup10 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    -- shared load operator group (11) : ptr_deref_2010_load_0 ptr_deref_2129_load_0 ptr_deref_2522_load_0 
    LoadGroup11: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2010_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2129_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2522_load_0_req_0;
      ptr_deref_2010_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2129_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2522_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2010_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2129_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2522_load_0_req_1;
      ptr_deref_2010_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2129_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2522_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup11_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup11_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup11_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup11_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup11_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup11_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup11_gI: SplitGuardInterface generic map(name => "LoadGroup11_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2010_word_address_0 & ptr_deref_2129_word_address_0 & ptr_deref_2522_word_address_0;
      ptr_deref_2010_data_0 <= data_out(95 downto 64);
      ptr_deref_2129_data_0 <= data_out(63 downto 32);
      ptr_deref_2522_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup11", addr_width => 10,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(9 downto 0),
          mtag => memory_space_1_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup11 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 11
    -- shared store operator group (0) : STORE_Nitr_required_2608_store_0 STORE_Nitr_required_2066_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_Nitr_required_2608_store_0_req_0;
      reqL_unguarded(0) <= STORE_Nitr_required_2066_store_0_req_0;
      STORE_Nitr_required_2608_store_0_ack_0 <= ackL_unguarded(1);
      STORE_Nitr_required_2066_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_Nitr_required_2608_store_0_req_1;
      reqR_unguarded(0) <= STORE_Nitr_required_2066_store_0_req_1;
      STORE_Nitr_required_2608_store_0_ack_1 <= ackR_unguarded(1);
      STORE_Nitr_required_2066_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_Nitr_required_2608_word_address_0 & STORE_Nitr_required_2066_word_address_0;
      data_in <= STORE_Nitr_required_2608_data_0 & STORE_Nitr_required_2066_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(15 downto 0),
          mtag => memory_space_0_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_is_decoded_2041_store_0 STORE_is_decoded_2169_store_0 STORE_is_decoded_2224_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= STORE_is_decoded_2041_store_0_req_0;
      reqL_unguarded(1) <= STORE_is_decoded_2169_store_0_req_0;
      reqL_unguarded(0) <= STORE_is_decoded_2224_store_0_req_0;
      STORE_is_decoded_2041_store_0_ack_0 <= ackL_unguarded(2);
      STORE_is_decoded_2169_store_0_ack_0 <= ackL_unguarded(1);
      STORE_is_decoded_2224_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= STORE_is_decoded_2041_store_0_req_1;
      reqR_unguarded(1) <= STORE_is_decoded_2169_store_0_req_1;
      reqR_unguarded(0) <= STORE_is_decoded_2224_store_0_req_1;
      STORE_is_decoded_2041_store_0_ack_1 <= ackR_unguarded(2);
      STORE_is_decoded_2169_store_0_ack_1 <= ackR_unguarded(1);
      STORE_is_decoded_2224_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_is_decoded_2041_word_address_0 & STORE_is_decoded_2169_word_address_0 & STORE_is_decoded_2224_word_address_0;
      data_in <= STORE_is_decoded_2041_data_0 & STORE_is_decoded_2169_data_0 & STORE_is_decoded_2224_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 0,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_2184_store_0 ptr_deref_1414_store_0 ptr_deref_2239_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 2, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 4, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2184_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1414_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2239_store_0_req_0;
      ptr_deref_2184_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1414_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2239_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2184_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1414_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2239_store_0_req_1;
      ptr_deref_2184_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1414_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2239_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2184_word_address_0 & ptr_deref_1414_word_address_0 & ptr_deref_2239_word_address_0;
      data_in <= ptr_deref_2184_data_0 & ptr_deref_1414_data_0 & ptr_deref_2239_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(9 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1538_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1538_store_0_req_0;
      ptr_deref_1538_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1538_store_0_req_1;
      ptr_deref_1538_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1538_word_address_0;
      data_in <= ptr_deref_1538_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(9 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_1667_store_0 ptr_deref_2544_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(19 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1667_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2544_store_0_req_0;
      ptr_deref_1667_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2544_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1667_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2544_store_0_req_1;
      ptr_deref_1667_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2544_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1667_word_address_0 & ptr_deref_2544_word_address_0;
      data_in <= ptr_deref_1667_data_0 & ptr_deref_2544_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(9 downto 0),
          mdata => memory_space_9_sr_data(31 downto 0),
          mtag => memory_space_9_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_2018_store_0 ptr_deref_1808_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(19 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2018_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1808_store_0_req_0;
      ptr_deref_2018_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1808_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2018_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1808_store_0_req_1;
      ptr_deref_2018_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1808_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2018_word_address_0 & ptr_deref_1808_word_address_0;
      data_in <= ptr_deref_2018_data_0 & ptr_deref_1808_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(9 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_1889_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1889_store_0_req_0;
      ptr_deref_1889_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1889_store_0_req_1;
      ptr_deref_1889_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1889_word_address_0;
      data_in <= ptr_deref_1889_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 10,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(9 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_code_block_in_1402_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_code_block_in_1402_inst_req_0;
      RPIPE_code_block_in_1402_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_code_block_in_1402_inst_req_1;
      RPIPE_code_block_in_1402_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iNsTr_17_1403 <= data_out(31 downto 0);
      code_block_in_read_0_gI: SplitGuardInterface generic map(name => "code_block_in_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      code_block_in_read_0: InputPortRevised -- 
        generic map ( name => "code_block_in_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => code_block_in_pipe_read_req(0),
          oack => code_block_in_pipe_read_ack(0),
          odata => code_block_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_code_block_decoded_2659_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_code_block_decoded_2659_inst_req_0;
      WPIPE_code_block_decoded_2659_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_code_block_decoded_2659_inst_req_1;
      WPIPE_code_block_decoded_2659_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= iNsTr_74_2658;
      code_block_decoded_write_0_gI: SplitGuardInterface generic map(name => "code_block_decoded_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      code_block_decoded_write_0: OutputPortRevised -- 
        generic map ( name => "code_block_decoded", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => code_block_decoded_pipe_write_req(0),
          oack => code_block_decoded_pipe_write_ack(0),
          odata => code_block_decoded_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nitr_required_2698_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nitr_required_2698_inst_req_0;
      WPIPE_nitr_required_2698_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nitr_required_2698_inst_req_1;
      WPIPE_nitr_required_2698_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= iNsTr_55_2689;
      nitr_required_write_1_gI: SplitGuardInterface generic map(name => "nitr_required_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nitr_required_write_1: OutputPortRevised -- 
        generic map ( name => "nitr_required", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nitr_required_pipe_write_req(0),
          oack => nitr_required_pipe_write_ack(0),
          odata => nitr_required_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1356_call 
    initInputs_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1356_call_req_0;
      call_stmt_1356_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1356_call_req_1;
      call_stmt_1356_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initInputs_call_group_0_gI: SplitGuardInterface generic map(name => "initInputs_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => initInputs_call_reqs(0),
          ackR => initInputs_call_acks(0),
          tagR => initInputs_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => initInputs_return_acks(0), -- cross-over
          ackL => initInputs_return_reqs(0), -- cross-over
          tagL => initInputs_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1913_call 
    checkNodeComputeEngine_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1913_call_req_0;
      call_stmt_1913_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1913_call_req_1;
      call_stmt_1913_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      checkNodeComputeEngine_call_group_1_gI: SplitGuardInterface generic map(name => "checkNodeComputeEngine_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => checkNodeComputeEngine_call_reqs(0),
          ackR => checkNodeComputeEngine_call_acks(0),
          tagR => checkNodeComputeEngine_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => checkNodeComputeEngine_return_acks(0), -- cross-over
          ackL => checkNodeComputeEngine_return_reqs(0), -- cross-over
          tagL => checkNodeComputeEngine_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end minSumDecode_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    code_block_decoded_pipe_read_data: out std_logic_vector(31 downto 0);
    code_block_decoded_pipe_read_req : in std_logic_vector(0 downto 0);
    code_block_decoded_pipe_read_ack : out std_logic_vector(0 downto 0);
    code_block_in_pipe_write_data: in std_logic_vector(31 downto 0);
    code_block_in_pipe_write_req : in std_logic_vector(0 downto 0);
    code_block_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_write_data: in std_logic_vector(31 downto 0);
    ebbyNo_in_pipe_write_req : in std_logic_vector(0 downto 0);
    ebbyNo_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    matrix_in_pipe_write_data: in std_logic_vector(15 downto 0);
    matrix_in_pipe_write_req : in std_logic_vector(0 downto 0);
    matrix_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxNitr_in_pipe_write_data: in std_logic_vector(15 downto 0);
    maxNitr_in_pipe_write_req : in std_logic_vector(0 downto 0);
    maxNitr_in_pipe_write_ack : out std_logic_vector(0 downto 0);
    nitr_required_pipe_read_data: out std_logic_vector(15 downto 0);
    nitr_required_pipe_read_req : in std_logic_vector(0 downto 0);
    nitr_required_pipe_read_ack : out std_logic_vector(0 downto 0);
    rate_in_pipe_write_data: in std_logic_vector(31 downto 0);
    rate_in_pipe_write_req : in std_logic_vector(0 downto 0);
    rate_in_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_10
  signal memory_space_10_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_10_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_10_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_10_lr_tag : std_logic_vector(9 downto 0);
  signal memory_space_10_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_10_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_10_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_10_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_11
  signal memory_space_11_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_11_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_11_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_12
  signal memory_space_12_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_12_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_12_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_12_lr_tag : std_logic_vector(9 downto 0);
  signal memory_space_12_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_12_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_12_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_12_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_12_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_12_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_12_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_13
  signal memory_space_13_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_13_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_13_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_13_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_13_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(19 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(9 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(29 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(47 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(8 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_9
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(9 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module checkNodeComputeEngine
  component checkNodeComputeEngine is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_9_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_9_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_9_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_9_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_12_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_12_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_12_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module checkNodeComputeEngine
  signal checkNodeComputeEngine_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal checkNodeComputeEngine_tag_out   : std_logic_vector(1 downto 0);
  signal checkNodeComputeEngine_start_req : std_logic;
  signal checkNodeComputeEngine_start_ack : std_logic;
  signal checkNodeComputeEngine_fin_req   : std_logic;
  signal checkNodeComputeEngine_fin_ack : std_logic;
  -- caller side aggregated signals for module checkNodeComputeEngine
  signal checkNodeComputeEngine_call_reqs: std_logic_vector(0 downto 0);
  signal checkNodeComputeEngine_call_acks: std_logic_vector(0 downto 0);
  signal checkNodeComputeEngine_return_reqs: std_logic_vector(0 downto 0);
  signal checkNodeComputeEngine_return_acks: std_logic_vector(0 downto 0);
  signal checkNodeComputeEngine_call_tag: std_logic_vector(0 downto 0);
  signal checkNodeComputeEngine_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module initInputs
  component initInputs is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_11_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_12_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_12_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_12_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_12_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_13_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_13_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_13_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_13_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_13_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_sc_tag :  in  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ebbyNo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      matrix_in_pipe_read_req : out  std_logic_vector(1 downto 0);
      matrix_in_pipe_read_ack : in   std_logic_vector(1 downto 0);
      matrix_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      maxNitr_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxNitr_in_pipe_read_data : in   std_logic_vector(15 downto 0);
      rate_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      rate_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rate_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initInputs
  signal initInputs_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initInputs_tag_out   : std_logic_vector(1 downto 0);
  signal initInputs_start_req : std_logic;
  signal initInputs_start_ack : std_logic;
  signal initInputs_fin_req   : std_logic;
  signal initInputs_fin_ack : std_logic;
  -- caller side aggregated signals for module initInputs
  signal initInputs_call_reqs: std_logic_vector(0 downto 0);
  signal initInputs_call_acks: std_logic_vector(0 downto 0);
  signal initInputs_return_reqs: std_logic_vector(0 downto 0);
  signal initInputs_return_acks: std_logic_vector(0 downto 0);
  signal initInputs_call_tag: std_logic_vector(0 downto 0);
  signal initInputs_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module minSumDecode
  component minSumDecode is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_11_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_11_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_11_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_11_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_11_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_11_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(9 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_12_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_12_lr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_12_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_12_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_12_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_12_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_13_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_13_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_13_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_13_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_13_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_13_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_13_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_9_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_9_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(5 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      code_block_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      code_block_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      code_block_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      code_block_decoded_pipe_write_req : out  std_logic_vector(0 downto 0);
      code_block_decoded_pipe_write_ack : in   std_logic_vector(0 downto 0);
      code_block_decoded_pipe_write_data : out  std_logic_vector(31 downto 0);
      nitr_required_pipe_write_req : out  std_logic_vector(0 downto 0);
      nitr_required_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nitr_required_pipe_write_data : out  std_logic_vector(15 downto 0);
      checkNodeComputeEngine_call_reqs : out  std_logic_vector(0 downto 0);
      checkNodeComputeEngine_call_acks : in   std_logic_vector(0 downto 0);
      checkNodeComputeEngine_call_tag  :  out  std_logic_vector(0 downto 0);
      checkNodeComputeEngine_return_reqs : out  std_logic_vector(0 downto 0);
      checkNodeComputeEngine_return_acks : in   std_logic_vector(0 downto 0);
      checkNodeComputeEngine_return_tag :  in   std_logic_vector(0 downto 0);
      initInputs_call_reqs : out  std_logic_vector(0 downto 0);
      initInputs_call_acks : in   std_logic_vector(0 downto 0);
      initInputs_call_tag  :  out  std_logic_vector(0 downto 0);
      initInputs_return_reqs : out  std_logic_vector(0 downto 0);
      initInputs_return_acks : in   std_logic_vector(0 downto 0);
      initInputs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module minSumDecode
  signal minSumDecode_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal minSumDecode_tag_out   : std_logic_vector(1 downto 0);
  signal minSumDecode_start_req : std_logic;
  signal minSumDecode_start_ack : std_logic;
  signal minSumDecode_fin_req   : std_logic;
  signal minSumDecode_fin_ack : std_logic;
  -- aggregate signals for write to pipe code_block_decoded
  signal code_block_decoded_pipe_write_data: std_logic_vector(31 downto 0);
  signal code_block_decoded_pipe_write_req: std_logic_vector(0 downto 0);
  signal code_block_decoded_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe code_block_in
  signal code_block_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal code_block_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal code_block_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ebbyNo_in
  signal ebbyNo_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal ebbyNo_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal ebbyNo_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe matrix_in
  signal matrix_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal matrix_in_pipe_read_req: std_logic_vector(1 downto 0);
  signal matrix_in_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe maxNitr_in
  signal maxNitr_in_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxNitr_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxNitr_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nitr_required
  signal nitr_required_pipe_write_data: std_logic_vector(15 downto 0);
  signal nitr_required_pipe_write_req: std_logic_vector(0 downto 0);
  signal nitr_required_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe rate_in
  signal rate_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal rate_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal rate_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module checkNodeComputeEngine
  -- call arbiter for module checkNodeComputeEngine
  checkNodeComputeEngine_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => checkNodeComputeEngine_call_reqs,
      call_acks => checkNodeComputeEngine_call_acks,
      return_reqs => checkNodeComputeEngine_return_reqs,
      return_acks => checkNodeComputeEngine_return_acks,
      call_tag  => checkNodeComputeEngine_call_tag,
      return_tag  => checkNodeComputeEngine_return_tag,
      call_mtag => checkNodeComputeEngine_tag_in,
      return_mtag => checkNodeComputeEngine_tag_out,
      call_mreq => checkNodeComputeEngine_start_req,
      call_mack => checkNodeComputeEngine_start_ack,
      return_mreq => checkNodeComputeEngine_fin_req,
      return_mack => checkNodeComputeEngine_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  checkNodeComputeEngine_instance:checkNodeComputeEngine-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => checkNodeComputeEngine_start_req,
      start_ack => checkNodeComputeEngine_start_ack,
      fin_req => checkNodeComputeEngine_fin_req,
      fin_ack => checkNodeComputeEngine_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_lr_req => memory_space_8_lr_req(2 downto 2),
      memory_space_8_lr_ack => memory_space_8_lr_ack(2 downto 2),
      memory_space_8_lr_addr => memory_space_8_lr_addr(29 downto 20),
      memory_space_8_lr_tag => memory_space_8_lr_tag(20 downto 14),
      memory_space_8_lc_req => memory_space_8_lc_req(2 downto 2),
      memory_space_8_lc_ack => memory_space_8_lc_ack(2 downto 2),
      memory_space_8_lc_data => memory_space_8_lc_data(47 downto 32),
      memory_space_8_lc_tag => memory_space_8_lc_tag(8 downto 6),
      memory_space_9_lr_req => memory_space_9_lr_req(0 downto 0),
      memory_space_9_lr_ack => memory_space_9_lr_ack(0 downto 0),
      memory_space_9_lr_addr => memory_space_9_lr_addr(9 downto 0),
      memory_space_9_lr_tag => memory_space_9_lr_tag(4 downto 0),
      memory_space_9_lc_req => memory_space_9_lc_req(0 downto 0),
      memory_space_9_lc_ack => memory_space_9_lc_ack(0 downto 0),
      memory_space_9_lc_data => memory_space_9_lc_data(31 downto 0),
      memory_space_9_lc_tag => memory_space_9_lc_tag(1 downto 0),
      memory_space_10_lr_req => memory_space_10_lr_req(1 downto 1),
      memory_space_10_lr_ack => memory_space_10_lr_ack(1 downto 1),
      memory_space_10_lr_addr => memory_space_10_lr_addr(1 downto 1),
      memory_space_10_lr_tag => memory_space_10_lr_tag(9 downto 5),
      memory_space_10_lc_req => memory_space_10_lc_req(1 downto 1),
      memory_space_10_lc_ack => memory_space_10_lc_ack(1 downto 1),
      memory_space_10_lc_data => memory_space_10_lc_data(31 downto 16),
      memory_space_10_lc_tag => memory_space_10_lc_tag(3 downto 2),
      memory_space_12_lr_req => memory_space_12_lr_req(1 downto 1),
      memory_space_12_lr_ack => memory_space_12_lr_ack(1 downto 1),
      memory_space_12_lr_addr => memory_space_12_lr_addr(1 downto 1),
      memory_space_12_lr_tag => memory_space_12_lr_tag(9 downto 5),
      memory_space_12_lc_req => memory_space_12_lc_req(1 downto 1),
      memory_space_12_lc_ack => memory_space_12_lc_ack(1 downto 1),
      memory_space_12_lc_data => memory_space_12_lc_data(31 downto 16),
      memory_space_12_lc_tag => memory_space_12_lc_tag(3 downto 2),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(19 downto 10),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 32),
      memory_space_5_sr_tag => memory_space_5_sr_tag(9 downto 5),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 2),
      tag_in => checkNodeComputeEngine_tag_in,
      tag_out => checkNodeComputeEngine_tag_out-- 
    ); -- 
  -- module initInputs
  -- call arbiter for module initInputs
  initInputs_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initInputs_call_reqs,
      call_acks => initInputs_call_acks,
      return_reqs => initInputs_return_reqs,
      return_acks => initInputs_return_acks,
      call_tag  => initInputs_call_tag,
      return_tag  => initInputs_return_tag,
      call_mtag => initInputs_tag_in,
      return_mtag => initInputs_tag_out,
      call_mreq => initInputs_start_req,
      call_mack => initInputs_start_ack,
      return_mreq => initInputs_fin_req,
      return_mack => initInputs_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  initInputs_instance:initInputs-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => initInputs_start_req,
      start_ack => initInputs_start_ack,
      fin_req => initInputs_fin_req,
      fin_ack => initInputs_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_lr_req => memory_space_8_lr_req(1 downto 1),
      memory_space_8_lr_ack => memory_space_8_lr_ack(1 downto 1),
      memory_space_8_lr_addr => memory_space_8_lr_addr(19 downto 10),
      memory_space_8_lr_tag => memory_space_8_lr_tag(13 downto 7),
      memory_space_8_lc_req => memory_space_8_lc_req(1 downto 1),
      memory_space_8_lc_ack => memory_space_8_lc_ack(1 downto 1),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 16),
      memory_space_8_lc_tag => memory_space_8_lc_tag(5 downto 3),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(3 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(3 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(9 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(6 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(2 downto 0),
      memory_space_10_sr_req => memory_space_10_sr_req(0 downto 0),
      memory_space_10_sr_ack => memory_space_10_sr_ack(0 downto 0),
      memory_space_10_sr_addr => memory_space_10_sr_addr(0 downto 0),
      memory_space_10_sr_data => memory_space_10_sr_data(15 downto 0),
      memory_space_10_sr_tag => memory_space_10_sr_tag(4 downto 0),
      memory_space_10_sc_req => memory_space_10_sc_req(0 downto 0),
      memory_space_10_sc_ack => memory_space_10_sc_ack(0 downto 0),
      memory_space_10_sc_tag => memory_space_10_sc_tag(1 downto 0),
      memory_space_11_sr_req => memory_space_11_sr_req(0 downto 0),
      memory_space_11_sr_ack => memory_space_11_sr_ack(0 downto 0),
      memory_space_11_sr_addr => memory_space_11_sr_addr(0 downto 0),
      memory_space_11_sr_data => memory_space_11_sr_data(15 downto 0),
      memory_space_11_sr_tag => memory_space_11_sr_tag(5 downto 0),
      memory_space_11_sc_req => memory_space_11_sc_req(0 downto 0),
      memory_space_11_sc_ack => memory_space_11_sc_ack(0 downto 0),
      memory_space_11_sc_tag => memory_space_11_sc_tag(2 downto 0),
      memory_space_12_sr_req => memory_space_12_sr_req(0 downto 0),
      memory_space_12_sr_ack => memory_space_12_sr_ack(0 downto 0),
      memory_space_12_sr_addr => memory_space_12_sr_addr(0 downto 0),
      memory_space_12_sr_data => memory_space_12_sr_data(15 downto 0),
      memory_space_12_sr_tag => memory_space_12_sr_tag(4 downto 0),
      memory_space_12_sc_req => memory_space_12_sc_req(0 downto 0),
      memory_space_12_sc_ack => memory_space_12_sc_ack(0 downto 0),
      memory_space_12_sc_tag => memory_space_12_sc_tag(1 downto 0),
      memory_space_13_sr_req => memory_space_13_sr_req(0 downto 0),
      memory_space_13_sr_ack => memory_space_13_sr_ack(0 downto 0),
      memory_space_13_sr_addr => memory_space_13_sr_addr(0 downto 0),
      memory_space_13_sr_data => memory_space_13_sr_data(31 downto 0),
      memory_space_13_sr_tag => memory_space_13_sr_tag(3 downto 0),
      memory_space_13_sc_req => memory_space_13_sc_req(0 downto 0),
      memory_space_13_sc_ack => memory_space_13_sc_ack(0 downto 0),
      memory_space_13_sc_tag => memory_space_13_sc_tag(0 downto 0),
      ebbyNo_in_pipe_read_req => ebbyNo_in_pipe_read_req(0 downto 0),
      ebbyNo_in_pipe_read_ack => ebbyNo_in_pipe_read_ack(0 downto 0),
      ebbyNo_in_pipe_read_data => ebbyNo_in_pipe_read_data(31 downto 0),
      matrix_in_pipe_read_req => matrix_in_pipe_read_req(1 downto 0),
      matrix_in_pipe_read_ack => matrix_in_pipe_read_ack(1 downto 0),
      matrix_in_pipe_read_data => matrix_in_pipe_read_data(31 downto 0),
      maxNitr_in_pipe_read_req => maxNitr_in_pipe_read_req(0 downto 0),
      maxNitr_in_pipe_read_ack => maxNitr_in_pipe_read_ack(0 downto 0),
      maxNitr_in_pipe_read_data => maxNitr_in_pipe_read_data(15 downto 0),
      rate_in_pipe_read_req => rate_in_pipe_read_req(0 downto 0),
      rate_in_pipe_read_ack => rate_in_pipe_read_ack(0 downto 0),
      rate_in_pipe_read_data => rate_in_pipe_read_data(31 downto 0),
      tag_in => initInputs_tag_in,
      tag_out => initInputs_tag_out-- 
    ); -- 
  -- module minSumDecode
  minSumDecode_instance:minSumDecode-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => minSumDecode_start_req,
      start_ack => minSumDecode_start_ack,
      fin_req => minSumDecode_fin_req,
      fin_ack => minSumDecode_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(4 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(15 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(9 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(4 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(9 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(4 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(9 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(5 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(3 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(9 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(4 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(1 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(3 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(9 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(6 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(15 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(2 downto 0),
      memory_space_10_lr_req => memory_space_10_lr_req(0 downto 0),
      memory_space_10_lr_ack => memory_space_10_lr_ack(0 downto 0),
      memory_space_10_lr_addr => memory_space_10_lr_addr(0 downto 0),
      memory_space_10_lr_tag => memory_space_10_lr_tag(4 downto 0),
      memory_space_10_lc_req => memory_space_10_lc_req(0 downto 0),
      memory_space_10_lc_ack => memory_space_10_lc_ack(0 downto 0),
      memory_space_10_lc_data => memory_space_10_lc_data(15 downto 0),
      memory_space_10_lc_tag => memory_space_10_lc_tag(1 downto 0),
      memory_space_11_lr_req => memory_space_11_lr_req(0 downto 0),
      memory_space_11_lr_ack => memory_space_11_lr_ack(0 downto 0),
      memory_space_11_lr_addr => memory_space_11_lr_addr(0 downto 0),
      memory_space_11_lr_tag => memory_space_11_lr_tag(5 downto 0),
      memory_space_11_lc_req => memory_space_11_lc_req(0 downto 0),
      memory_space_11_lc_ack => memory_space_11_lc_ack(0 downto 0),
      memory_space_11_lc_data => memory_space_11_lc_data(15 downto 0),
      memory_space_11_lc_tag => memory_space_11_lc_tag(2 downto 0),
      memory_space_12_lr_req => memory_space_12_lr_req(0 downto 0),
      memory_space_12_lr_ack => memory_space_12_lr_ack(0 downto 0),
      memory_space_12_lr_addr => memory_space_12_lr_addr(0 downto 0),
      memory_space_12_lr_tag => memory_space_12_lr_tag(4 downto 0),
      memory_space_12_lc_req => memory_space_12_lc_req(0 downto 0),
      memory_space_12_lc_ack => memory_space_12_lc_ack(0 downto 0),
      memory_space_12_lc_data => memory_space_12_lc_data(15 downto 0),
      memory_space_12_lc_tag => memory_space_12_lc_tag(1 downto 0),
      memory_space_13_lr_req => memory_space_13_lr_req(0 downto 0),
      memory_space_13_lr_ack => memory_space_13_lr_ack(0 downto 0),
      memory_space_13_lr_addr => memory_space_13_lr_addr(0 downto 0),
      memory_space_13_lr_tag => memory_space_13_lr_tag(3 downto 0),
      memory_space_13_lc_req => memory_space_13_lc_req(0 downto 0),
      memory_space_13_lc_ack => memory_space_13_lc_ack(0 downto 0),
      memory_space_13_lc_data => memory_space_13_lc_data(31 downto 0),
      memory_space_13_lc_tag => memory_space_13_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(15 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(4 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(9 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(4 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(9 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(4 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(9 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(5 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(9 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(4 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(1 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 0),
      memory_space_9_sr_req => memory_space_9_sr_req(0 downto 0),
      memory_space_9_sr_ack => memory_space_9_sr_ack(0 downto 0),
      memory_space_9_sr_addr => memory_space_9_sr_addr(9 downto 0),
      memory_space_9_sr_data => memory_space_9_sr_data(31 downto 0),
      memory_space_9_sr_tag => memory_space_9_sr_tag(4 downto 0),
      memory_space_9_sc_req => memory_space_9_sc_req(0 downto 0),
      memory_space_9_sc_ack => memory_space_9_sc_ack(0 downto 0),
      memory_space_9_sc_tag => memory_space_9_sc_tag(1 downto 0),
      code_block_in_pipe_read_req => code_block_in_pipe_read_req(0 downto 0),
      code_block_in_pipe_read_ack => code_block_in_pipe_read_ack(0 downto 0),
      code_block_in_pipe_read_data => code_block_in_pipe_read_data(31 downto 0),
      code_block_decoded_pipe_write_req => code_block_decoded_pipe_write_req(0 downto 0),
      code_block_decoded_pipe_write_ack => code_block_decoded_pipe_write_ack(0 downto 0),
      code_block_decoded_pipe_write_data => code_block_decoded_pipe_write_data(31 downto 0),
      nitr_required_pipe_write_req => nitr_required_pipe_write_req(0 downto 0),
      nitr_required_pipe_write_ack => nitr_required_pipe_write_ack(0 downto 0),
      nitr_required_pipe_write_data => nitr_required_pipe_write_data(15 downto 0),
      checkNodeComputeEngine_call_reqs => checkNodeComputeEngine_call_reqs(0 downto 0),
      checkNodeComputeEngine_call_acks => checkNodeComputeEngine_call_acks(0 downto 0),
      checkNodeComputeEngine_call_tag => checkNodeComputeEngine_call_tag(0 downto 0),
      checkNodeComputeEngine_return_reqs => checkNodeComputeEngine_return_reqs(0 downto 0),
      checkNodeComputeEngine_return_acks => checkNodeComputeEngine_return_acks(0 downto 0),
      checkNodeComputeEngine_return_tag => checkNodeComputeEngine_return_tag(0 downto 0),
      initInputs_call_reqs => initInputs_call_reqs(0 downto 0),
      initInputs_call_acks => initInputs_call_acks(0 downto 0),
      initInputs_call_tag => initInputs_call_tag(0 downto 0),
      initInputs_return_reqs => initInputs_return_reqs(0 downto 0),
      initInputs_return_acks => initInputs_return_acks(0 downto 0),
      initInputs_return_tag => initInputs_return_tag(0 downto 0),
      tag_in => minSumDecode_tag_in,
      tag_out => minSumDecode_tag_out-- 
    ); -- 
  -- module will be run forever 
  minSumDecode_tag_in <= (others => '0');
  minSumDecode_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => minSumDecode_start_req, start_ack => minSumDecode_start_ack,  fin_req => minSumDecode_fin_req,  fin_ack => minSumDecode_fin_ack);
  code_block_decoded_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe code_block_decoded",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => code_block_decoded_pipe_read_req,
      read_ack => code_block_decoded_pipe_read_ack,
      read_data => code_block_decoded_pipe_read_data,
      write_req => code_block_decoded_pipe_write_req,
      write_ack => code_block_decoded_pipe_write_ack,
      write_data => code_block_decoded_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  code_block_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe code_block_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => code_block_in_pipe_read_req,
      read_ack => code_block_in_pipe_read_ack,
      read_data => code_block_in_pipe_read_data,
      write_req => code_block_in_pipe_write_req,
      write_ack => code_block_in_pipe_write_ack,
      write_data => code_block_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ebbyNo_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ebbyNo_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => ebbyNo_in_pipe_read_req,
      read_ack => ebbyNo_in_pipe_read_ack,
      read_data => ebbyNo_in_pipe_read_data,
      write_req => ebbyNo_in_pipe_write_req,
      write_ack => ebbyNo_in_pipe_write_ack,
      write_data => ebbyNo_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  matrix_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe matrix_in",
      num_reads => 2,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => matrix_in_pipe_read_req,
      read_ack => matrix_in_pipe_read_ack,
      read_data => matrix_in_pipe_read_data,
      write_req => matrix_in_pipe_write_req,
      write_ack => matrix_in_pipe_write_ack,
      write_data => matrix_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxNitr_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxNitr_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxNitr_in_pipe_read_req,
      read_ack => maxNitr_in_pipe_read_ack,
      read_data => maxNitr_in_pipe_read_data,
      write_req => maxNitr_in_pipe_write_req,
      write_ack => maxNitr_in_pipe_write_ack,
      write_data => maxNitr_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nitr_required_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nitr_required",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => nitr_required_pipe_read_req,
      read_ack => nitr_required_pipe_read_ack,
      read_data => nitr_required_pipe_read_data,
      write_req => nitr_required_pipe_write_req,
      write_ack => nitr_required_pipe_write_ack,
      write_data => nitr_required_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  rate_in_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe rate_in",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      depth => 2 --
    )
    port map( -- 
      read_req => rate_in_pipe_read_req,
      read_ack => rate_in_pipe_read_ack,
      read_data => rate_in_pipe_read_data,
      write_req => rate_in_pipe_write_req,
      write_ack => rate_in_pipe_write_ack,
      write_data => rate_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_10: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_10",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_10_lr_addr,
      lr_req_in => memory_space_10_lr_req,
      lr_ack_out => memory_space_10_lr_ack,
      lr_tag_in => memory_space_10_lr_tag,
      lc_req_in => memory_space_10_lc_req,
      lc_ack_out => memory_space_10_lc_ack,
      lc_data_out => memory_space_10_lc_data,
      lc_tag_out => memory_space_10_lc_tag,
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_11: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_11",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_11_lr_addr,
      lr_req_in => memory_space_11_lr_req,
      lr_ack_out => memory_space_11_lr_ack,
      lr_tag_in => memory_space_11_lr_tag,
      lc_req_in => memory_space_11_lc_req,
      lc_ack_out => memory_space_11_lc_ack,
      lc_data_out => memory_space_11_lc_data,
      lc_tag_out => memory_space_11_lc_tag,
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_12: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_12",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_12_lr_addr,
      lr_req_in => memory_space_12_lr_req,
      lr_ack_out => memory_space_12_lr_ack,
      lr_tag_in => memory_space_12_lr_tag,
      lc_req_in => memory_space_12_lc_req,
      lc_ack_out => memory_space_12_lc_ack,
      lc_data_out => memory_space_12_lc_data,
      lc_tag_out => memory_space_12_lc_tag,
      sr_addr_in => memory_space_12_sr_addr,
      sr_data_in => memory_space_12_sr_data,
      sr_req_in => memory_space_12_sr_req,
      sr_ack_out => memory_space_12_sr_ack,
      sr_tag_in => memory_space_12_sr_tag,
      sc_req_in=> memory_space_12_sc_req,
      sc_ack_out => memory_space_12_sc_ack,
      sc_tag_out => memory_space_12_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_13: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_13",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_13_lr_addr,
      lr_req_in => memory_space_13_lr_req,
      lr_ack_out => memory_space_13_lr_ack,
      lr_tag_in => memory_space_13_lr_tag,
      lc_req_in => memory_space_13_lc_req,
      lc_ack_out => memory_space_13_lc_ack,
      lc_data_out => memory_space_13_lc_data,
      lc_tag_out => memory_space_13_lc_tag,
      sr_addr_in => memory_space_13_sr_addr,
      sr_data_in => memory_space_13_sr_data,
      sr_req_in => memory_space_13_sr_req,
      sr_ack_out => memory_space_13_sr_ack,
      sr_tag_in => memory_space_13_sr_tag,
      sc_req_in=> memory_space_13_sc_req,
      sc_ack_out => memory_space_13_sc_ack,
      sc_tag_out => memory_space_13_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 2,
      addr_width => 10,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_6: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 3,
      num_stores => 1,
      addr_width => 10,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 4,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_9",
      num_loads => 1,
      num_stores => 1,
      addr_width => 10,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 10,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
