-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant Nitr_required_base_address : std_logic_vector(0 downto 0) := "0";
  constant aPosteriori_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant aPriori_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant code_block_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant ebbyNo_base_address : std_logic_vector(0 downto 0) := "0";
  constant ext_info_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant is_decoded_base_address : std_logic_vector(0 downto 0) := "0";
  constant maxNitr_base_address : std_logic_vector(0 downto 0) := "0";
  constant mem_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant message_base_address : std_logic_vector(9 downto 0) := "0000000000";
  constant ncol_ind_base_address : std_logic_vector(0 downto 0) := "0";
  constant ncols_base_address : std_logic_vector(0 downto 0) := "0";
  constant nrows_base_address : std_logic_vector(0 downto 0) := "0";
  constant rate_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package ahir_system_global_package;
